`timescale 1ns/1ps
`default_nettype wire
module fe65p2 ( I2536792601E6CADEAB49502F1BD19044 , IB5859D8721CFDC0312B2838B9C985BC1
,I0657423B4C5BA1BD8F1054E02912833A , IB8CD801B107A9A8F62C5B61EA5646620 , I816D49F5014DFDC552FDCBE11E19B458 , I236DDEB5A953C3C3F6AC87852A12F153 , I1BAD808A5C69D4BE6F74A54F1DB10784 ,
I97EB8C7F0ADCF2A52AECB93D7E606AD4 , I8CCA42A31A8386AF5CCBA8CAE1E7580B , I1F5748542B5178997408DBA54D0F2CD3 , ICC25F554E80352BF341B28E9BA1E817F ,
I38CB737AD9DAD35E6421516AE85D9130 , I13A780F88690EA17740517649EB0E7C5 , I6CC01EBE09C98E8D2223196A8E4D7A6A , IC00738DF0D4BEC8A1C8ED0B3ABAB3881 , IF962DDDFCFB59F7648E592F6EAE19C93 ,
I0ED2ADDC6F83E144925F05986E9CFF86 , IA95AE92E4828AF7B0DADD49D537FEE5E , I958F38294CE0C6337C616E28CE0C0EF4 , I531D5C1FBCF6E356CAFEEBA55A5B73D0 ,
I3405A5272BCD250BE6AAB2071FA8E2C7 , I0F71A3473EE22B4B3DACA05365112EB4 , IE3B0A4C4EA55DD2B44B6B72D7B0966A2 , I2F93BC5D4AA9CC738D29F51E46D80581 ,
I6F8FB1BAF897A3508E8CE28CC0047AFE , I5E982716C925AA53DFAD54323E066CD2 , I154AA2DDCB3DAA94E8CBB3AC8C7CB247 , I5B9F987DBE3EDAC4E347A14A5782131F ,
I08C038534302D663980480E37D20BC83 , I769454D2A8D191F3E322B7B5DF928B5D , I01BDC194686F6DC3F502CFA733822312 , I87B3D78A5F6FFC46951ED28E772E594D ,
I159859469876028CEA112C7C16B1CAF5 , IAE766072895E2EB8B8716944E133AE63 ); input wire [64*64-1:0] I2536792601E6CADEAB49502F1BD19044 ; input
wire [1:0] IB5859D8721CFDC0312B2838B9C985BC1 ; input wire I0657423B4C5BA1BD8F1054E02912833A , IB8CD801B107A9A8F62C5B61EA5646620 ; input
wire I1BAD808A5C69D4BE6F74A54F1DB10784 , I97EB8C7F0ADCF2A52AECB93D7E606AD4 , I8CCA42A31A8386AF5CCBA8CAE1E7580B ,
I1F5748542B5178997408DBA54D0F2CD3 ; output reg ICC25F554E80352BF341B28E9BA1E817F ; input wire I13A780F88690EA17740517649EB0E7C5 ; output
wire I6CC01EBE09C98E8D2223196A8E4D7A6A , IC00738DF0D4BEC8A1C8ED0B3ABAB3881 ; input wire I38CB737AD9DAD35E6421516AE85D9130 ; output
wire I816D49F5014DFDC552FDCBE11E19B458 , I236DDEB5A953C3C3F6AC87852A12F153 ; input wire IF962DDDFCFB59F7648E592F6EAE19C93 ;
inout wire I0ED2ADDC6F83E144925F05986E9CFF86 , IA95AE92E4828AF7B0DADD49D537FEE5E , I958F38294CE0C6337C616E28CE0C0EF4 ,
I531D5C1FBCF6E356CAFEEBA55A5B73D0 , I3405A5272BCD250BE6AAB2071FA8E2C7 , I0F71A3473EE22B4B3DACA05365112EB4 , IE3B0A4C4EA55DD2B44B6B72D7B0966A2 ,
I2F93BC5D4AA9CC738D29F51E46D80581 , I6F8FB1BAF897A3508E8CE28CC0047AFE , I5E982716C925AA53DFAD54323E066CD2 , I154AA2DDCB3DAA94E8CBB3AC8C7CB247 ; localparam
I54C65A028FF224383655ADAB430D6741 = 16; inout wire [I54C65A028FF224383655ADAB430D6741 *2-1:0] I5B9F987DBE3EDAC4E347A14A5782131F ,
I08C038534302D663980480E37D20BC83 , I769454D2A8D191F3E322B7B5DF928B5D , I01BDC194686F6DC3F502CFA733822312 , I87B3D78A5F6FFC46951ED28E772E594D ,
I159859469876028CEA112C7C16B1CAF5 ; output wire [63:0] IAE766072895E2EB8B8716944E133AE63 ; wire IF37891DFD06D53B7D2C58D80CE50E1EC ; wire
I4032B1FC75E1EC6D7B4EC5F598A8CCA8 ; assign I816D49F5014DFDC552FDCBE11E19B458 = IF37891DFD06D53B7D2C58D80CE50E1EC ; assign
I236DDEB5A953C3C3F6AC87852A12F153 = !IF37891DFD06D53B7D2C58D80CE50E1EC ; assign I6CC01EBE09C98E8D2223196A8E4D7A6A
= I4032B1FC75E1EC6D7B4EC5F598A8CCA8 ; assign IC00738DF0D4BEC8A1C8ED0B3ABAB3881 = !I4032B1FC75E1EC6D7B4EC5F598A8CCA8 ; reg
IAEA9A05B5360FCBA85A008A029FFD1E2 ; wire I361CDAC76AF22A4F90CFCDB9BC018036 ; reg I92A3CB8DEDEC0EBEE60321250DF1BB8A ; reg
I435F5BE3A446834FFCDFBF8C61E7B715 ; wire I3309F577FB69AF63D0F9276438540F1F ; reg I3D22F82428FBB3DDBC3F1007022E8882 ; reg
I6990F9296B2B9B77E498A7417648BDD7 ; reg I06081CF6EEC3FACFA54ED9EC41EC568A ; always @(*) begin if (I97EB8C7F0ADCF2A52AECB93D7E606AD4 )
begin I3D22F82428FBB3DDBC3F1007022E8882 = I1F5748542B5178997408DBA54D0F2CD3 ; I6990F9296B2B9B77E498A7417648BDD7
= I8CCA42A31A8386AF5CCBA8CAE1E7580B ; I06081CF6EEC3FACFA54ED9EC41EC568A = I1BAD808A5C69D4BE6F74A54F1DB10784 ; IAEA9A05B5360FCBA85A008A029FFD1E2
= 0; I92A3CB8DEDEC0EBEE60321250DF1BB8A = 0; I435F5BE3A446834FFCDFBF8C61E7B715 = 0; ICC25F554E80352BF341B28E9BA1E817F
= I3309F577FB69AF63D0F9276438540F1F ; end else begin I3D22F82428FBB3DDBC3F1007022E8882 = 0; I6990F9296B2B9B77E498A7417648BDD7
= 0; I06081CF6EEC3FACFA54ED9EC41EC568A = 0; IAEA9A05B5360FCBA85A008A029FFD1E2 = I1F5748542B5178997408DBA54D0F2CD3 ; I92A3CB8DEDEC0EBEE60321250DF1BB8A
= I8CCA42A31A8386AF5CCBA8CAE1E7580B ; I435F5BE3A446834FFCDFBF8C61E7B715 = I1BAD808A5C69D4BE6F74A54F1DB10784 ; ICC25F554E80352BF341B28E9BA1E817F
= I361CDAC76AF22A4F90CFCDB9BC018036 ; end end reg ID31AA1C2707092E408AE9E599CC3A844 , I8EB85E51C21BED1CE594F9D9162709AA ,
I1A5D8348640CD64ABC78C0F8236DE0D5 ; always @(*) begin if (IB5859D8721CFDC0312B2838B9C985BC1 == 2'b00) begin ID31AA1C2707092E408AE9E599CC3A844
= 0; I8EB85E51C21BED1CE594F9D9162709AA = 1; I1A5D8348640CD64ABC78C0F8236DE0D5 = 1; end else if (IB5859D8721CFDC0312B2838B9C985BC1
== 2'b01) begin ID31AA1C2707092E408AE9E599CC3A844 = 1; I8EB85E51C21BED1CE594F9D9162709AA = 0; I1A5D8348640CD64ABC78C0F8236DE0D5
= 0; end else if (IB5859D8721CFDC0312B2838B9C985BC1 == 2'b10) begin ID31AA1C2707092E408AE9E599CC3A844 = 0; I8EB85E51C21BED1CE594F9D9162709AA
= 1; I1A5D8348640CD64ABC78C0F8236DE0D5 = 0; end else begin ID31AA1C2707092E408AE9E599CC3A844 = 0; I8EB85E51C21BED1CE594F9D9162709AA
= 0; I1A5D8348640CD64ABC78C0F8236DE0D5 = 0; end end localparam I7AAD85FA8F0E841E1283EBD8BA7E3285 = 145; wire [I7AAD85FA8F0E841E1283EBD8BA7E3285 -1:0]
I59041103AA4B47824D6D362D800C06DA , IB9E9A17061E48936432FE29691D71CEE , I89A166B2AF2BC9835FD1510FB08C5273 ; I9BBBBEA9F740C6E76E42F55F5AB2A5A2
#(.I62E5CEF85D46F1A5A2144D9FD463B79E (I7AAD85FA8F0E841E1283EBD8BA7E3285 )) I0467BCB3142906DD43F3481C41AE850F ( .I0EB8CC186C9B38B7FB99E477EE981265 (I8EB85E51C21BED1CE594F9D9162709AA ),
.I0A3BC2148686F2B562665C3891507E35 (I435F5BE3A446834FFCDFBF8C61E7B715 ), .I946490AD0FDC17B3B899760A445128F0 (I92A3CB8DEDEC0EBEE60321250DF1BB8A ),
.IAC5585D98646D255299C359140537783 (IAEA9A05B5360FCBA85A008A029FFD1E2 ), .IB807023F87E63B8ADA92F79F546FF9CC (I361CDAC76AF22A4F90CFCDB9BC018036 ), .I08804A5B28516A9DC9E56ABFEECF66D9 (I59041103AA4B47824D6D362D800C06DA ),
.I7C147CDA9E49590F6ABE83D118B7353B (IB9E9A17061E48936432FE29691D71CEE ), .IE78AFF6FF490ECAC5AFE4B8DF2BDC999 (I89A166B2AF2BC9835FD1510FB08C5273 ) ); wire
I102B0AB51A9FDD94E90B3701B6BE31CE ; wire I6742A038F36525E7B03E8A1E9E5FEDB4 ; wire ID3D904FD6B5F5F28BE04E2A4E0A7E103 ; wire
[3:0] I2812F2D69AFEDB8661D5EC3468BF8B29 ; wire [1:0] I54D5B5297D6861DCB70E3BC023CF557D ; wire [1:0] I8357B924AEFCA0FDD29AADC1ABE078FF ; wire
[8:0] I22C3EC380D38314B0801D994F39EF010 ; wire [15:0] I3F9C583C4A9E941ACBE85A2594F7E352 ; wire [15:0] ICE93BBB963818B0EF722D742F12E5637 ; wire
[3:0] I018E74A6510FFC837EA6A71BA2E4CB09 ; wire I1C95AC4E3DEEA066549E9C90BCB0C1E0 ; wire [7:0] I11F95A0C5F7742674A79BC87E1B2964D ,
I84084D39F62AE5D8A52B11B1253ABCDE , I162409FF040F7F3E2DA52B937D494D30 , ID3A582311A8E071B679C274DBDFD7215 , I5C233C51F04AD0630FF42B367E8683C0 ,
I6984213466AAA84C606C16C53C3E605A , I2BE6E12A300F68CF67FEF00D8AA324B9 , IF67A010C8FC31412C9C71C06D18C03F1 , IA630490703D6C7FC3EA60013645C6089 ,
I7C6A8ECC7AB01190AB26356C01FE1D2C , I06A4C8E444893BE261332501F9CEDF79 ; assign I102B0AB51A9FDD94E90B3701B6BE31CE
= I89A166B2AF2BC9835FD1510FB08C5273 [0]; assign I6742A038F36525E7B03E8A1E9E5FEDB4 = I89A166B2AF2BC9835FD1510FB08C5273 [1]; assign
ID3D904FD6B5F5F28BE04E2A4E0A7E103 = I89A166B2AF2BC9835FD1510FB08C5273 [2]; assign I2812F2D69AFEDB8661D5EC3468BF8B29
= I89A166B2AF2BC9835FD1510FB08C5273 [6:3]; assign I54D5B5297D6861DCB70E3BC023CF557D = I89A166B2AF2BC9835FD1510FB08C5273 [8:7]; assign
I1C95AC4E3DEEA066549E9C90BCB0C1E0 = IB9E9A17061E48936432FE29691D71CEE [10]; assign I59041103AA4B47824D6D362D800C06DA [10]
= 1; assign I22C3EC380D38314B0801D994F39EF010 = IB9E9A17061E48936432FE29691D71CEE [20:12]; assign I59041103AA4B47824D6D362D800C06DA [20:12]
= 401; assign I3F9C583C4A9E941ACBE85A2594F7E352 = IB9E9A17061E48936432FE29691D71CEE [36:21]; assign I59041103AA4B47824D6D362D800C06DA [36:21]
= 16'hffff; assign ICE93BBB963818B0EF722D742F12E5637 = IB9E9A17061E48936432FE29691D71CEE [52:37]; assign I59041103AA4B47824D6D362D800C06DA [52:37]
= 16'hffff; assign I018E74A6510FFC837EA6A71BA2E4CB09 = IB9E9A17061E48936432FE29691D71CEE [56:53]; assign I59041103AA4B47824D6D362D800C06DA [56:53]
= 15; assign I11F95A0C5F7742674A79BC87E1B2964D = IB9E9A17061E48936432FE29691D71CEE [64:57]; assign I59041103AA4B47824D6D362D800C06DA [64:57]
= 0; assign I84084D39F62AE5D8A52B11B1253ABCDE = IB9E9A17061E48936432FE29691D71CEE [72:65]; assign I59041103AA4B47824D6D362D800C06DA [72:65]
= 36; assign I162409FF040F7F3E2DA52B937D494D30 = IB9E9A17061E48936432FE29691D71CEE [80:73]; assign I59041103AA4B47824D6D362D800C06DA [80:73]
= 255; assign ID3A582311A8E071B679C274DBDFD7215 = IB9E9A17061E48936432FE29691D71CEE [88:81]; assign I59041103AA4B47824D6D362D800C06DA [88:81]
= 0; assign I5C233C51F04AD0630FF42B367E8683C0 = IB9E9A17061E48936432FE29691D71CEE [96:89]; assign I59041103AA4B47824D6D362D800C06DA [96:89]
= 42; assign I6984213466AAA84C606C16C53C3E605A = IB9E9A17061E48936432FE29691D71CEE [104:97]; assign I59041103AA4B47824D6D362D800C06DA [104:97]
= 0; assign I2BE6E12A300F68CF67FEF00D8AA324B9 = IB9E9A17061E48936432FE29691D71CEE [112:105]; assign I59041103AA4B47824D6D362D800C06DA [112:105]
= 0; assign IF67A010C8FC31412C9C71C06D18C03F1 = IB9E9A17061E48936432FE29691D71CEE [120:113]; assign I59041103AA4B47824D6D362D800C06DA [120:113]
= 51; assign IA630490703D6C7FC3EA60013645C6089 = IB9E9A17061E48936432FE29691D71CEE [128:121]; assign I59041103AA4B47824D6D362D800C06DA [128:121]
= 1; assign I7C6A8ECC7AB01190AB26356C01FE1D2C = IB9E9A17061E48936432FE29691D71CEE [136:129]; assign I59041103AA4B47824D6D362D800C06DA [136:129]
= 25; assign I06A4C8E444893BE261332501F9CEDF79 = IB9E9A17061E48936432FE29691D71CEE [144:137]; assign I59041103AA4B47824D6D362D800C06DA [144:137]
= 50; wire I21345BCEA5A3A0213882E3493F7CE8A2 , IE8F9438C61FEFC48890126E846737803 , I00D170E901FDFA8C4D428ECAC839A4AB ; wire
[3:0] I182E80B21C5A5F086FE70D9A01554365 ; wire [1:0] I453DD3088EE862556BDD0F58B390F41F ; assign I21345BCEA5A3A0213882E3493F7CE8A2
= I102B0AB51A9FDD94E90B3701B6BE31CE & I92A3CB8DEDEC0EBEE60321250DF1BB8A ; assign IE8F9438C61FEFC48890126E846737803
= I6742A038F36525E7B03E8A1E9E5FEDB4 & I92A3CB8DEDEC0EBEE60321250DF1BB8A ; assign I00D170E901FDFA8C4D428ECAC839A4AB
= ID3D904FD6B5F5F28BE04E2A4E0A7E103 & I92A3CB8DEDEC0EBEE60321250DF1BB8A ; assign I182E80B21C5A5F086FE70D9A01554365
= I2812F2D69AFEDB8661D5EC3468BF8B29 & {4{I92A3CB8DEDEC0EBEE60321250DF1BB8A }}; assign I453DD3088EE862556BDD0F58B390F41F
= I54D5B5297D6861DCB70E3BC023CF557D & {2{I92A3CB8DEDEC0EBEE60321250DF1BB8A }}; wire [1:0] I9B7ED19526E1EF8476E81C4995389C4D ,
I696DE38724D3F45226B3BFADCA2221B0 , I2942DAE8F4C3E4D7DE62D00DF109B597 , IBD4BC8D76A5E12444220433B31B0D5AE , I4E230A7B3BA8125AC46C2C29E4ED732C ,
I862FFD9F0CD7DD281B24BCD321EF5998 , I3270527819CE05DB94D853B81288E61E , I7F429D68386CA0F2B2233B532306EAFA , IA775ECF21554187489A5ADE053F04828 ,
IDDA1F0A1D5E5A6BB9E09B84272ED69B9 , IF4090A076C6B2B05DFED25AD11AA6619 ; assign I0ED2ADDC6F83E144925F05986E9CFF86
= |I84084D39F62AE5D8A52B11B1253ABCDE ; assign IA95AE92E4828AF7B0DADD49D537FEE5E = |I162409FF040F7F3E2DA52B937D494D30 ; assign
I958F38294CE0C6337C616E28CE0C0EF4 = |ID3A582311A8E071B679C274DBDFD7215 ; assign I531D5C1FBCF6E356CAFEEBA55A5B73D0
= |I5C233C51F04AD0630FF42B367E8683C0 ; assign I3405A5272BCD250BE6AAB2071FA8E2C7 = |I6984213466AAA84C606C16C53C3E605A ; assign
I0F71A3473EE22B4B3DACA05365112EB4 = |I2BE6E12A300F68CF67FEF00D8AA324B9 ; assign IE3B0A4C4EA55DD2B44B6B72D7B0966A2
= |IF67A010C8FC31412C9C71C06D18C03F1 ; assign I2F93BC5D4AA9CC738D29F51E46D80581 = |IA630490703D6C7FC3EA60013645C6089 ; assign
I6F8FB1BAF897A3508E8CE28CC0047AFE = |I7C6A8ECC7AB01190AB26356C01FE1D2C ; assign I5E982716C925AA53DFAD54323E066CD2
= |I06A4C8E444893BE261332501F9CEDF79 ; assign I9B7ED19526E1EF8476E81C4995389C4D = {2{IF962DDDFCFB59F7648E592F6EAE19C93 }}; assign
I696DE38724D3F45226B3BFADCA2221B0 = {2{I0ED2ADDC6F83E144925F05986E9CFF86 }}; assign I2942DAE8F4C3E4D7DE62D00DF109B597
= {2{IA95AE92E4828AF7B0DADD49D537FEE5E }}; assign IBD4BC8D76A5E12444220433B31B0D5AE = {2{I958F38294CE0C6337C616E28CE0C0EF4 }}; assign
I4E230A7B3BA8125AC46C2C29E4ED732C = {2{I531D5C1FBCF6E356CAFEEBA55A5B73D0 }}; assign I862FFD9F0CD7DD281B24BCD321EF5998
= {2{I3405A5272BCD250BE6AAB2071FA8E2C7 }}; assign I3270527819CE05DB94D853B81288E61E = {2{I0F71A3473EE22B4B3DACA05365112EB4 }}; assign
I7F429D68386CA0F2B2233B532306EAFA = {2{IE3B0A4C4EA55DD2B44B6B72D7B0966A2 }}; assign IA775ECF21554187489A5ADE053F04828
= {2{I2F93BC5D4AA9CC738D29F51E46D80581 }}; assign IDDA1F0A1D5E5A6BB9E09B84272ED69B9 = {2{I6F8FB1BAF897A3508E8CE28CC0047AFE }}; assign
IF4090A076C6B2B05DFED25AD11AA6619 = {2{I5E982716C925AA53DFAD54323E066CD2 }}; wire [15:0] IF6068DAA29DBB05A7EAD1E3B5A48BBEE ; wire
[5:0] IA70367AA7CB74E510F4F9413CCF059D3 ; wire [3:0] I1976D7F704DE389D9FE064E08EA35B2D ; wire [15:0] IB69F2E4AAFE438766DDFFC3511700FCB
[I54C65A028FF224383655ADAB430D6741 -1:0]; wire [5:0] IF5A84EE8549E66B9C336DCF93F594D98 [I54C65A028FF224383655ADAB430D6741 -1:0]; assign
IF6068DAA29DBB05A7EAD1E3B5A48BBEE = IB69F2E4AAFE438766DDFFC3511700FCB [0] | IB69F2E4AAFE438766DDFFC3511700FCB [1]
| IB69F2E4AAFE438766DDFFC3511700FCB [2] | IB69F2E4AAFE438766DDFFC3511700FCB [3] | IB69F2E4AAFE438766DDFFC3511700FCB [4]
| IB69F2E4AAFE438766DDFFC3511700FCB [5] | IB69F2E4AAFE438766DDFFC3511700FCB [6] | IB69F2E4AAFE438766DDFFC3511700FCB [7]
| IB69F2E4AAFE438766DDFFC3511700FCB [8] | IB69F2E4AAFE438766DDFFC3511700FCB [9] | IB69F2E4AAFE438766DDFFC3511700FCB [10]
| IB69F2E4AAFE438766DDFFC3511700FCB [11] | IB69F2E4AAFE438766DDFFC3511700FCB [12] | IB69F2E4AAFE438766DDFFC3511700FCB [13]
| IB69F2E4AAFE438766DDFFC3511700FCB [14] | IB69F2E4AAFE438766DDFFC3511700FCB [15] ; assign IA70367AA7CB74E510F4F9413CCF059D3
= IF5A84EE8549E66B9C336DCF93F594D98 [0] | IF5A84EE8549E66B9C336DCF93F594D98 [1] | IF5A84EE8549E66B9C336DCF93F594D98 [2]
| IF5A84EE8549E66B9C336DCF93F594D98 [3] | IF5A84EE8549E66B9C336DCF93F594D98 [4] | IF5A84EE8549E66B9C336DCF93F594D98 [5]
| IF5A84EE8549E66B9C336DCF93F594D98 [6] | IF5A84EE8549E66B9C336DCF93F594D98 [7] | IF5A84EE8549E66B9C336DCF93F594D98 [8]
| IF5A84EE8549E66B9C336DCF93F594D98 [9] | IF5A84EE8549E66B9C336DCF93F594D98 [10] | IF5A84EE8549E66B9C336DCF93F594D98 [11]
| IF5A84EE8549E66B9C336DCF93F594D98 [12] | IF5A84EE8549E66B9C336DCF93F594D98 [13] | IF5A84EE8549E66B9C336DCF93F594D98 [14]
| IF5A84EE8549E66B9C336DCF93F594D98 [15] ; wire [3:0] I0590CD3F1ABD6DC5F1FAF1EE1CB75731 [I54C65A028FF224383655ADAB430D6741 :0]; assign
I0590CD3F1ABD6DC5F1FAF1EE1CB75731 [0] = 0; assign I1976D7F704DE389D9FE064E08EA35B2D = I0590CD3F1ABD6DC5F1FAF1EE1CB75731 [I54C65A028FF224383655ADAB430D6741 ]; wire
I94A08DA1FECBB6E8B46990538C7B50B2 ; wire [I54C65A028FF224383655ADAB430D6741 :0] IA2C5BD9372B8600132A16A5093637C36 ; assign
IA2C5BD9372B8600132A16A5093637C36 [0] = 0; assign I94A08DA1FECBB6E8B46990538C7B50B2 = IA2C5BD9372B8600132A16A5093637C36 [I54C65A028FF224383655ADAB430D6741 ]; wire
[I54C65A028FF224383655ADAB430D6741 -1:0] I804B8A3C0F4E36EB8002981FA0CC4F12 ; assign I3309F577FB69AF63D0F9276438540F1F
= I804B8A3C0F4E36EB8002981FA0CC4F12 [I018E74A6510FFC837EA6A71BA2E4CB09 ]; wire [I54C65A028FF224383655ADAB430D6741 -1:0]
I48A355561F0628CB2813BD54EADAA46C , I64C0936E5F806DE5E4330429CC8ACC6D ; assign I64C0936E5F806DE5E4330429CC8ACC6D
= I48A355561F0628CB2813BD54EADAA46C & I3F9C583C4A9E941ACBE85A2594F7E352 ; assign IF37891DFD06D53B7D2C58D80CE50E1EC
= |I64C0936E5F806DE5E4330429CC8ACC6D ; wire IC3C311DE1CD01CDF3D31BB00F2B0E9E2 ; wire IEDB112AE72B861E77CF4D55A756C76FC ; wire
[3:0] IE9DED2DF97E91174FD62E40E248B137D , I8715FEDE1A202C700CD025C90F3B2421 ; reg [8:0] I082A499B7DDEF3C7897AB842B431A8AD ,
I89C5B8F33C91378743762C771A89F8C4 ; reg [I54C65A028FF224383655ADAB430D6741 -1:0] I02A145553791DED7486E3D55412998B3 ; always @(*)
begin if (I1C95AC4E3DEEA066549E9C90BCB0C1E0 ) I02A145553791DED7486E3D55412998B3 = {I804B8A3C0F4E36EB8002981FA0CC4F12 [I54C65A028FF224383655ADAB430D6741 -2:0],
I3D22F82428FBB3DDBC3F1007022E8882 }; else I02A145553791DED7486E3D55412998B3 = ICE93BBB963818B0EF722D742F12E5637
& {16{I3D22F82428FBB3DDBC3F1007022E8882 }}; end `ifndef TEST_DC
localparam I24140871F9CD6D3D93FBAAB2DB509EBB = I54C65A028FF224383655ADAB430D6741 ; `else
localparam I24140871F9CD6D3D93FBAAB2DB509EBB = `TEST_DC;
`endif
wire [63:0] I5367F16813E8B3314F5C3786E492456F [I54C65A028FF224383655ADAB430D6741 -1:0]; assign IAE766072895E2EB8B8716944E133AE63
= I5367F16813E8B3314F5C3786E492456F [I54C65A028FF224383655ADAB430D6741 -1]; generate genvar I8CE4B16B22B58894AA86C421E8759DF3 ; for
(I8CE4B16B22B58894AA86C421E8759DF3 =0; I8CE4B16B22B58894AA86C421E8759DF3 <I54C65A028FF224383655ADAB430D6741 ; I8CE4B16B22B58894AA86C421E8759DF3 =I8CE4B16B22B58894AA86C421E8759DF3 +1) begin :
IE689416A84F62A67F362E7C637AC05F8 wire IE2E897D79A478206E8991CE3054B1B01 = I3F9C583C4A9E941ACBE85A2594F7E352 [I8CE4B16B22B58894AA86C421E8759DF3 ]; wire
I199366DFFA7738F8028B2DD0CA3E78A0 = ICE93BBB963818B0EF722D742F12E5637 [I8CE4B16B22B58894AA86C421E8759DF3 ]; wire
IAE23F82FE849CA57AFF8C2B976AB930E ; wire ID09326563FB1E5A3A6598AAF65A746C2 ; wire [15:0] I0EF1C97DC12E8501873AFD9288FB4F66 ; wire
[5:0] I1BDFD64578BF098597347B27C098F615 ; assign IB69F2E4AAFE438766DDFFC3511700FCB [I8CE4B16B22B58894AA86C421E8759DF3 ]
= (IAE23F82FE849CA57AFF8C2B976AB930E & IE2E897D79A478206E8991CE3054B1B01 ) ? I0EF1C97DC12E8501873AFD9288FB4F66 :
0; assign IF5A84EE8549E66B9C336DCF93F594D98 [I8CE4B16B22B58894AA86C421E8759DF3 ] = (IAE23F82FE849CA57AFF8C2B976AB930E
& IE2E897D79A478206E8991CE3054B1B01 ) ? I1BDFD64578BF098597347B27C098F615 : 0; if (I8CE4B16B22B58894AA86C421E8759DF3
<I24140871F9CD6D3D93FBAAB2DB509EBB ) begin I21F5A4F10878160CE707AC6682B91D1B I5F11B53FF7202633EA278395908DB7DA ( .I2536792601E6CADEAB49502F1BD19044 (I2536792601E6CADEAB49502F1BD19044 [(I8CE4B16B22B58894AA86C421E8759DF3 +1)*(64*4)-1:I8CE4B16B22B58894AA86C421E8759DF3 *(64*4)]), .I27E9DD9482B253AA850544215471D9D5 (IC3C311DE1CD01CDF3D31BB00F2B0E9E2
& IE2E897D79A478206E8991CE3054B1B01 ), .I86266EE937D97F812A8E57D22B62EE29 (ID31AA1C2707092E408AE9E599CC3A844 ) ,.I0A3BC2148686F2B562665C3891507E35 (I0657423B4C5BA1BD8F1054E02912833A
& IE2E897D79A478206E8991CE3054B1B01 ), .I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 (IAE23F82FE849CA57AFF8C2B976AB930E & IE2E897D79A478206E8991CE3054B1B01 ),
.IE9DED2DF97E91174FD62E40E248B137D (IE9DED2DF97E91174FD62E40E248B137D & {4{IE2E897D79A478206E8991CE3054B1B01 }}),
.I8715FEDE1A202C700CD025C90F3B2421 (I8715FEDE1A202C700CD025C90F3B2421 & {4{IE2E897D79A478206E8991CE3054B1B01 }}),
.I1A7B4E094F07B0C85C5ACADEC807841F (ID09326563FB1E5A3A6598AAF65A746C2 ), .I21345BCEA5A3A0213882E3493F7CE8A2 (I21345BCEA5A3A0213882E3493F7CE8A2
& I199366DFFA7738F8028B2DD0CA3E78A0 ), .IE8F9438C61FEFC48890126E846737803 (IE8F9438C61FEFC48890126E846737803 & I199366DFFA7738F8028B2DD0CA3E78A0 ),
.I00D170E901FDFA8C4D428ECAC839A4AB (I00D170E901FDFA8C4D428ECAC839A4AB & I199366DFFA7738F8028B2DD0CA3E78A0 ), .I453DD3088EE862556BDD0F58B390F41F (I453DD3088EE862556BDD0F58B390F41F
& {2{I199366DFFA7738F8028B2DD0CA3E78A0 }}), .I182E80B21C5A5F086FE70D9A01554365 (I182E80B21C5A5F086FE70D9A01554365
& {4{I199366DFFA7738F8028B2DD0CA3E78A0 }}), .I346A81471C889B6C72A88423EB28B21A (I38CB737AD9DAD35E6421516AE85D9130 ),
.I0EB8CC186C9B38B7FB99E477EE981265 (I1A5D8348640CD64ABC78C0F8236DE0D5 ), .IF41F5F2D34464C2F1512CE4A38EAD286 (I06081CF6EEC3FACFA54ED9EC41EC568A
& I199366DFFA7738F8028B2DD0CA3E78A0 ), .I75D612F1AEBBE1DC3FC1AC2ED5C21E7F (I97EB8C7F0ADCF2A52AECB93D7E606AD4 & I199366DFFA7738F8028B2DD0CA3E78A0 ),
.IA882574F5206B0DBAB0B61BA8B369A15 (I02A145553791DED7486E3D55412998B3 [I8CE4B16B22B58894AA86C421E8759DF3 ]), .IE78AFF6FF490ECAC5AFE4B8DF2BDC999 (I804B8A3C0F4E36EB8002981FA0CC4F12 [I8CE4B16B22B58894AA86C421E8759DF3 ]),
.I24D24CDA7F2D8B539E4F5C420BD826D9 (I48A355561F0628CB2813BD54EADAA46C [I8CE4B16B22B58894AA86C421E8759DF3 ]), .I082A499B7DDEF3C7897AB842B431A8AD (I082A499B7DDEF3C7897AB842B431A8AD
& {9{IE2E897D79A478206E8991CE3054B1B01 }}), .I89C5B8F33C91378743762C771A89F8C4 (I89C5B8F33C91378743762C771A89F8C4
& {9{IE2E897D79A478206E8991CE3054B1B01 }}), .I8357B924AEFCA0FDD29AADC1ABE078FF (I8357B924AEFCA0FDD29AADC1ABE078FF ), .IF6068DAA29DBB05A7EAD1E3B5A48BBEE (I0EF1C97DC12E8501873AFD9288FB4F66 ),
.IA70367AA7CB74E510F4F9413CCF059D3 (I1BDFD64578BF098597347B27C098F615 ), .I61BAAAAF32AC5A7B6FFEBFC244A2D739 (I9B7ED19526E1EF8476E81C4995389C4D ),
.I6E03B4F12533CBA29903F1C9DD1E5C3D (I696DE38724D3F45226B3BFADCA2221B0 ), .IAB9D6A507309488CCF13DB3F67F81B63 (I2942DAE8F4C3E4D7DE62D00DF109B597 ),
.I83FCEFDFE9F9D1C28AB321626447799F (IBD4BC8D76A5E12444220433B31B0D5AE ), .I1905DD05FA116073F500B593198EED1C (I4E230A7B3BA8125AC46C2C29E4ED732C ),
.I61E6EBA71A6BFA5A8FE92AB8FABECBBC (I862FFD9F0CD7DD281B24BCD321EF5998 ), .I79EB40C7CC07F0A913BA2E8F9D56D33B (I3270527819CE05DB94D853B81288E61E ),
.I973092C325E8C2AE92FFF50B0288E777 (I7F429D68386CA0F2B2233B532306EAFA ), .IB9445BEC437AE377554E2723C22C52B2 (IA775ECF21554187489A5ADE053F04828 ),
.I6A45CBE320E935B06BB0F08ECF1179D4 (IDDA1F0A1D5E5A6BB9E09B84272ED69B9 ), .I0EE48206D3023D05A5AA46FD33711C98 (IF4090A076C6B2B05DFED25AD11AA6619 ), .I81414FA30C7BC73A9A778574097A714B (I9B7ED19526E1EF8476E81C4995389C4D ),
.I4C39D6D4449338A7DA014742DE16FD46 (I696DE38724D3F45226B3BFADCA2221B0 ), .ID8E8746A568679217650DF444D98F91E (I2942DAE8F4C3E4D7DE62D00DF109B597 ),
.I30CD5687FB19DAD9CFD43FE994021B00 (IBD4BC8D76A5E12444220433B31B0D5AE ), .I018477AF087A1484F83E54C386C2EF07 (I4E230A7B3BA8125AC46C2C29E4ED732C ),
.I6970ADE3C1C5CEF4BF2ADF425B8B73CB (I862FFD9F0CD7DD281B24BCD321EF5998 ), .I4021D2C4A029457D9671036AF92F0AB8 (I3270527819CE05DB94D853B81288E61E ),
.I6ABED3933223BDB35402C9F56973AB09 (I7F429D68386CA0F2B2233B532306EAFA ), .I371CC04BDE216A35CEFED5553951955B (IA775ECF21554187489A5ADE053F04828 ),
.I032B17AEE0B7BC21B073F5A5AF886D30 (IDDA1F0A1D5E5A6BB9E09B84272ED69B9 ), .I64571D3B8AD6548BEF3F326B0C79154D (IF4090A076C6B2B05DFED25AD11AA6619 ), .I5B9F987DBE3EDAC4E347A14A5782131F (I5B9F987DBE3EDAC4E347A14A5782131F [2*I8CE4B16B22B58894AA86C421E8759DF3 +1:2*I8CE4B16B22B58894AA86C421E8759DF3 ]),
.I08C038534302D663980480E37D20BC83 (I08C038534302D663980480E37D20BC83 [2*I8CE4B16B22B58894AA86C421E8759DF3 +1:2*I8CE4B16B22B58894AA86C421E8759DF3 ]), .I769454D2A8D191F3E322B7B5DF928B5D (I769454D2A8D191F3E322B7B5DF928B5D [2*I8CE4B16B22B58894AA86C421E8759DF3 +1:2*I8CE4B16B22B58894AA86C421E8759DF3 ]),
.I01BDC194686F6DC3F502CFA733822312 (I01BDC194686F6DC3F502CFA733822312 [2*I8CE4B16B22B58894AA86C421E8759DF3 +1:2*I8CE4B16B22B58894AA86C421E8759DF3 ]),
.I87B3D78A5F6FFC46951ED28E772E594D (I87B3D78A5F6FFC46951ED28E772E594D [2*I8CE4B16B22B58894AA86C421E8759DF3 +1:2*I8CE4B16B22B58894AA86C421E8759DF3 ]),
.I159859469876028CEA112C7C16B1CAF5 (I159859469876028CEA112C7C16B1CAF5 [2*I8CE4B16B22B58894AA86C421E8759DF3 +1:2*I8CE4B16B22B58894AA86C421E8759DF3 ]), .IAE766072895E2EB8B8716944E133AE63 (I5367F16813E8B3314F5C3786E492456F [I8CE4B16B22B58894AA86C421E8759DF3 ]) ); end else
begin assign ID09326563FB1E5A3A6598AAF65A746C2 = 0; end IFDB931B30D7BFF08B173BCF1F98E495C #(.I2664F03AC6B8BB9EEE4287720E407DB3 (I8CE4B16B22B58894AA86C421E8759DF3 ))
I670C28811C37FB7B943F1AEF363C9A49 ( .I586A6D64D60A5A9D3DD45E81AA6585A3 (IA2C5BD9372B8600132A16A5093637C36 [I8CE4B16B22B58894AA86C421E8759DF3 ]), .I2E192DB878F41E38E0F3B32CFC289D8F (ID09326563FB1E5A3A6598AAF65A746C2 ),
.I002953A92DEB31BDFD9E165DFB1DFE1C (IA2C5BD9372B8600132A16A5093637C36 [I8CE4B16B22B58894AA86C421E8759DF3 +1]), .I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 (IEDB112AE72B861E77CF4D55A756C76FC ),
.IAE23F82FE849CA57AFF8C2B976AB930E (IAE23F82FE849CA57AFF8C2B976AB930E ), .IA5CFBE42922BF86EC0D0DC539D627112 (I0590CD3F1ABD6DC5F1FAF1EE1CB75731 [I8CE4B16B22B58894AA86C421E8759DF3 +1]),
.IFA829BE14FC3FF9B411978DBF7DDF9EE (I0590CD3F1ABD6DC5F1FAF1EE1CB75731 [I8CE4B16B22B58894AA86C421E8759DF3 ]) ); end endgenerate reg
[8:0] IAD63AE7192A86A295FF0D6A7D7A79A67 ; wire [8:0] I18D3ECEEDB3A4C2EF443AFC3C82BC50A ; always @(posedge I0657423B4C5BA1BD8F1054E02912833A ) if (ID31AA1C2707092E408AE9E599CC3A844 ) IAD63AE7192A86A295FF0D6A7D7A79A67
<= 0; else IAD63AE7192A86A295FF0D6A7D7A79A67 <= IAD63AE7192A86A295FF0D6A7D7A79A67 + 1; assign I18D3ECEEDB3A4C2EF443AFC3C82BC50A
= IAD63AE7192A86A295FF0D6A7D7A79A67 - I22C3EC380D38314B0801D994F39EF010 ; always @(posedge I0657423B4C5BA1BD8F1054E02912833A ) #5ns
I082A499B7DDEF3C7897AB842B431A8AD <= (IAD63AE7192A86A295FF0D6A7D7A79A67 >> 1) ^ IAD63AE7192A86A295FF0D6A7D7A79A67 ; always @(posedge
I0657423B4C5BA1BD8F1054E02912833A ) #5ns I89C5B8F33C91378743762C771A89F8C4 <= (I18D3ECEEDB3A4C2EF443AFC3C82BC50A
>> 1) ^ I18D3ECEEDB3A4C2EF443AFC3C82BC50A ; wire I2320407509CCCBDA7D63F6D622F67DD8 , I38778258922E1E4431B75D526DC701D3 ;
wire [23:0] IE55603E44DA0CE59B3E8963A06AA6E5A ; wire ICB7658367C9FDD7110EBE09C34077D2C , I2AE05249E15E8C6BF7F6AB2A4306FACA ; reg
I9B343CDCB441F7E0267501DFEC7F7CBB ; I67D38CAA7C80960859CB2AFCF45A4106 I39EE20CB79819AB0991598E6D8FC4024 ( .I86266EE937D97F812A8E57D22B62EE29 (ID31AA1C2707092E408AE9E599CC3A844 ),
.I0A3BC2148686F2B562665C3891507E35 (I0657423B4C5BA1BD8F1054E02912833A ), .IF698F67F5666AFF10729D8A1CB1C14D2 (IB8CD801B107A9A8F62C5B61EA5646620 ),
.I459A6F79AD9B13CBCB5F692D2CC7A94D (I94A08DA1FECBB6E8B46990538C7B50B2 ), .IE7D31FC0602FB2EDE144D18CDFFD816B (!I38778258922E1E4431B75D526DC701D3
& !I9B343CDCB441F7E0267501DFEC7F7CBB ), .I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 (IEDB112AE72B861E77CF4D55A756C76FC ),
.I2C0F741D5E54A03052A7BAEB8CEFA690 (IC3C311DE1CD01CDF3D31BB00F2B0E9E2 ), .I43938353D4FB12C9720D1A7A7537E069 (IE9DED2DF97E91174FD62E40E248B137D ),
.I6413911CE482DB3AB245D5F066541602 (I8715FEDE1A202C700CD025C90F3B2421 ), .IE55603E44DA0CE59B3E8963A06AA6E5A (IE55603E44DA0CE59B3E8963A06AA6E5A ), .ICB7658367C9FDD7110EBE09C34077D2C (ICB7658367C9FDD7110EBE09C34077D2C ),
.I2AE05249E15E8C6BF7F6AB2A4306FACA (I2AE05249E15E8C6BF7F6AB2A4306FACA ), .IC68AD92486D949E2FF7EE4E70CD71E8E () ); reg
[25:0] IEB020EACC0DB5519E339450779B0AF6B ; wire [25:0] I9448935ECF6E007795136E89B711630A ; reg [25:0] I4BFA1D1EE173176C7AF5C2500CE29F70 ; wire
[3:0] I1A2BF9DFB7CD7E97B9849E2F2C053E63 [3:0]; assign I1A2BF9DFB7CD7E97B9849E2F2C053E63 [3] = IF6068DAA29DBB05A7EAD1E3B5A48BBEE [15:12]; assign
I1A2BF9DFB7CD7E97B9849E2F2C053E63 [2] = IF6068DAA29DBB05A7EAD1E3B5A48BBEE [11:8]; assign I1A2BF9DFB7CD7E97B9849E2F2C053E63 [1]
= IF6068DAA29DBB05A7EAD1E3B5A48BBEE [7:4]; assign I1A2BF9DFB7CD7E97B9849E2F2C053E63 [0] = IF6068DAA29DBB05A7EAD1E3B5A48BBEE [3:0]; assign
I9448935ECF6E007795136E89B711630A = {1'b0, 1'b0, 1'b0, 2'b0, I1976D7F704DE389D9FE064E08EA35B2D [3:0], IA70367AA7CB74E510F4F9413CCF059D3 [5:0],
1'b0, 2'b0, I1A2BF9DFB7CD7E97B9849E2F2C053E63 [3], I1A2BF9DFB7CD7E97B9849E2F2C053E63 [2]}; always @(posedge I0657423B4C5BA1BD8F1054E02912833A )
begin if (ICB7658367C9FDD7110EBE09C34077D2C ) I4BFA1D1EE173176C7AF5C2500CE29F70 <= {1'b0, 1'b0, 1'b0, 2'b0, I1976D7F704DE389D9FE064E08EA35B2D [3:0],
IA70367AA7CB74E510F4F9413CCF059D3 [5:0], 1'b1, 2'b0, I1A2BF9DFB7CD7E97B9849E2F2C053E63 [1], I1A2BF9DFB7CD7E97B9849E2F2C053E63 [0]}; end wire
I8F54A08C6D22B69A16FB31012E3B47A3 ; assign I8F54A08C6D22B69A16FB31012E3B47A3 = I2AE05249E15E8C6BF7F6AB2A4306FACA
| I9B343CDCB441F7E0267501DFEC7F7CBB | ICB7658367C9FDD7110EBE09C34077D2C ; always @(posedge I0657423B4C5BA1BD8F1054E02912833A )
begin if (ID31AA1C2707092E408AE9E599CC3A844 ) I9B343CDCB441F7E0267501DFEC7F7CBB <= 0; else if (ICB7658367C9FDD7110EBE09C34077D2C ) I9B343CDCB441F7E0267501DFEC7F7CBB
<= 1; else if (I9B343CDCB441F7E0267501DFEC7F7CBB & !I38778258922E1E4431B75D526DC701D3 ) I9B343CDCB441F7E0267501DFEC7F7CBB
<= 0; end always @(*) begin IEB020EACC0DB5519E339450779B0AF6B = 0; if (I2AE05249E15E8C6BF7F6AB2A4306FACA ) IEB020EACC0DB5519E339450779B0AF6B
= {1'b1,1'b0, 1'b1, IE55603E44DA0CE59B3E8963A06AA6E5A [22:0]}; if (ICB7658367C9FDD7110EBE09C34077D2C ) IEB020EACC0DB5519E339450779B0AF6B
= I9448935ECF6E007795136E89B711630A ; if (I9B343CDCB441F7E0267501DFEC7F7CBB ) IEB020EACC0DB5519E339450779B0AF6B
= I4BFA1D1EE173176C7AF5C2500CE29F70 ; end wire I5924C0A7318E32EE219C181624EDEA2D , IEA7B6999CAE148C37168B2D2F3EAC05B ,
IBD800844D88AC36F7C86D5A16D4BB69F ; wire [25:0] I93E489D255515612291AB619A9BC3041 ; reg [2:0] IBCD62779E44421FB36165DD34952DC2B ; always @(posedge
I0657423B4C5BA1BD8F1054E02912833A ) IBCD62779E44421FB36165DD34952DC2B <= {IBCD62779E44421FB36165DD34952DC2B [1:0],
ID31AA1C2707092E408AE9E599CC3A844 }; I4A7799F98F8BFA916086832ADA73E798 #(.I6DF7E246C71D6D2493823379E5C1AA50 (26),
.IDBF04E8E8F1F83557BAE7BEA2CBD57BD (3)) IA338F4828952E69A833F4AC5F8747427 ( .I5316F360783B270FE9AC3887CE27EF1D (I93E489D255515612291AB619A9BC3041 ), .IE01D0BDC7D5682BCB747F7EEFBE73DCB (I38778258922E1E4431B75D526DC701D3 ), .I561AF95BF4F6EB0D6654C5812AB28B1F (I5924C0A7318E32EE219C181624EDEA2D ), .IA776DD7EA52A4C6B834F3E481B7BDC1F (IEB020EACC0DB5519E339450779B0AF6B ), .I72A3034E1DBCB3283E6B3211A628FBD8 (I8F54A08C6D22B69A16FB31012E3B47A3 ),
.I9AB96B3F1E8B9326C3C792CB4B2BA759 (I0657423B4C5BA1BD8F1054E02912833A ), .I5814C91DB64F071BEEAA8913CE4B41D9 (ID31AA1C2707092E408AE9E599CC3A844 ), .I9B05D4C8F2C4E4DEE91A9C511A75634B (IEA7B6999CAE148C37168B2D2F3EAC05B ),
.I444A7039B02C6D02C8913AA00CF03207 (IBD800844D88AC36F7C86D5A16D4BB69F ), .I480B3FA2D679840798F74A04A6C7C705 (IBCD62779E44421FB36165DD34952DC2B [2]) ); wire
ID57871DE58E6EE367F695170D2090779 ; assign ID57871DE58E6EE367F695170D2090779 = I93E489D255515612291AB619A9BC3041 [25]; I507DE87DD0643D9F2D064D87FF8CE8DD
IBB1015E3BE27EBB1B06ECBA6E2258FAB ( .I86266EE937D97F812A8E57D22B62EE29 (ID31AA1C2707092E408AE9E599CC3A844 ), .I0A3BC2148686F2B562665C3891507E35 (I13A780F88690EA17740517649EB0E7C5 ),
.ID9C51D9F54B5E373B300DA2EDDDBB764 (I5924C0A7318E32EE219C181624EDEA2D ), .I8D777F385D3DFEC8815D20F7496026DC (I93E489D255515612291AB619A9BC3041 [23:0]), .I231E0CDCBF2977BEA26AECDA5A7F45FC (IEA7B6999CAE148C37168B2D2F3EAC05B ), .I3D2E8D60C335C528A7C12445BD1F41E3 (IBD800844D88AC36F7C86D5A16D4BB69F ), .IC68271A63DDBC431C307BEB7D2918275 (I4032B1FC75E1EC6D7B4EC5F598A8CCA8 ), .I50BB776CBF75FDBDD857EF107CDA97D3 (1'b0), .IB4702C9059470087164094C2E5F94070 (1'b0), .IA55086E1186D1C3CC0FFF510278DF91E (8'b0), .IB61F32A2FFDFF16751219654FC5AE6E7 (ID57871DE58E6EE367F695170D2090779 ) );
endmodule module IEF91D04B90E6EC355FF6DD49C50BA7EA (I7694F4A66316E53C8CDD9D9954BD611D , I0A3BC2148686F2B562665C3891507E35 ,
ICDAEEEBA9B4A4C5EBF042C0215A7BB0E ); output reg I7694F4A66316E53C8CDD9D9954BD611D ; input wire I0A3BC2148686F2B562665C3891507E35 ;
input wire ICDAEEEBA9B4A4C5EBF042C0215A7BB0E ; always @ (negedge I0A3BC2148686F2B562665C3891507E35 or posedge ICDAEEEBA9B4A4C5EBF042C0215A7BB0E ) if (ICDAEEEBA9B4A4C5EBF042C0215A7BB0E ) I7694F4A66316E53C8CDD9D9954BD611D
<= 1; else I7694F4A66316E53C8CDD9D9954BD611D <= !I7694F4A66316E53C8CDD9D9954BD611D ; endmodule module I6CCBE3F36B144174D7B5131F1612067F (IABEB1D6F727D4016CBA8D230E06173E2 ,
I975E762C6BF4B17F34E0966F54272008 , I37D350E5B2683ED4E78F696D8B080140 , ICFE6055D2E0503BE378BB63449EC7BA6 , IECAE13117D6F0584C25A9DA6C8F8415E ,
I8D777F385D3DFEC8815D20F7496026DC , I0A3BC2148686F2B562665C3891507E35 , I86266EE937D97F812A8E57D22B62EE29 , ID6299EFF2098B99E8BB408F652A2EE38 ,
I4CA8F5C40F80B904A3A115368EF165BF , I8357B924AEFCA0FDD29AADC1ABE078FF ); input wire IABEB1D6F727D4016CBA8D230E06173E2 ,
ICFE6055D2E0503BE378BB63449EC7BA6 , I0A3BC2148686F2B562665C3891507E35 , I86266EE937D97F812A8E57D22B62EE29 , ID6299EFF2098B99E8BB408F652A2EE38 ; output
wire I975E762C6BF4B17F34E0966F54272008 , I4CA8F5C40F80B904A3A115368EF165BF ; input wire [6:0] IECAE13117D6F0584C25A9DA6C8F8415E ; input
wire [6:0] I37D350E5B2683ED4E78F696D8B080140 ; output wire [3:0] I8D777F385D3DFEC8815D20F7496026DC ; input wire
[1:0] I8357B924AEFCA0FDD29AADC1ABE078FF ; wire [3:0] I288F847370AB993102C86AB98BD79E53 ; reg [2:0] I3776F996EEB88CF403041684C2E146BB ; wire
I7A640F52E5CF4CEF5E9DFB04D8BC271A ; assign I7A640F52E5CF4CEF5E9DFB04D8BC271A = IABEB1D6F727D4016CBA8D230E06173E2
| (|I3776F996EEB88CF403041684C2E146BB ) ; wire I8DE2A9CF71BCBDDB6996310B6090B645 ; I379BDABA1FBE95FD8A49051997E9665F
IF3A4CB21DB974338EEBF1A1CE7CFD675 (.I6F13D2E1112161FE6F8EA1EDD3F01310 (I0A3BC2148686F2B562665C3891507E35 ), .I208F156D4A803025C284BB595A7576B4 (I7A640F52E5CF4CEF5E9DFB04D8BC271A
| ICFE6055D2E0503BE378BB63449EC7BA6 ), .I3F3B6F139F935CDE0338584380A06130 (I8DE2A9CF71BCBDDB6996310B6090B645 )); always
@ (posedge I8DE2A9CF71BCBDDB6996310B6090B645 or posedge I86266EE937D97F812A8E57D22B62EE29 ) begin : ICD2ABC221E1D3CBABE06F94DFB93798A if (I86266EE937D97F812A8E57D22B62EE29 ) I3776F996EEB88CF403041684C2E146BB [2:0]
<= 0; else I3776F996EEB88CF403041684C2E146BB [2:0] <= { IABEB1D6F727D4016CBA8D230E06173E2 , I3776F996EEB88CF403041684C2E146BB [2:1]
}; end wire I76A88EC8C7A9140348BA5E2DAEEC0E89 ; assign I76A88EC8C7A9140348BA5E2DAEEC0E89 = I3776F996EEB88CF403041684C2E146BB [1:0]
== 2'b10; wire I0D28BD8A8650B66243673EBB8D515084 ; assign I0D28BD8A8650B66243673EBB8D515084 = I3776F996EEB88CF403041684C2E146BB [1:0]
== 2'b01; wire I25DC7640AC100AF468B94F57FF6E466A ; wire IB8B590EE84AE0766462AEF1DB7759CDF ; assign IB8B590EE84AE0766462AEF1DB7759CDF
= (I3776F996EEB88CF403041684C2E146BB [1] & !(I288F847370AB993102C86AB98BD79E53 == 4'd14)); I379BDABA1FBE95FD8A49051997E9665F
I0ADD073B14B25AF2A5E28C6D824C8D2E (.I6F13D2E1112161FE6F8EA1EDD3F01310 (I8DE2A9CF71BCBDDB6996310B6090B645 ), .I208F156D4A803025C284BB595A7576B4 (IB8B590EE84AE0766462AEF1DB7759CDF ),
.I3F3B6F139F935CDE0338584380A06130 (I25DC7640AC100AF468B94F57FF6E466A )); wire ID39228DB5F904D97CC6F69301B95F2D9 ; assign
ID39228DB5F904D97CC6F69301B95F2D9 = I86266EE937D97F812A8E57D22B62EE29 | (I3776F996EEB88CF403041684C2E146BB [2:1]
== 2'b10); IEF91D04B90E6EC355FF6DD49C50BA7EA I9F3FCC1B61D824135F8841AD9EF2A5BF (.I7694F4A66316E53C8CDD9D9954BD611D (I288F847370AB993102C86AB98BD79E53 [0]),
.I0A3BC2148686F2B562665C3891507E35 (I25DC7640AC100AF468B94F57FF6E466A ), .ICDAEEEBA9B4A4C5EBF042C0215A7BB0E (ID39228DB5F904D97CC6F69301B95F2D9 )); IEF91D04B90E6EC355FF6DD49C50BA7EA
I11EA41312F79DA5ADF9180387FEBBF73 (.I7694F4A66316E53C8CDD9D9954BD611D (I288F847370AB993102C86AB98BD79E53 [1]), .I0A3BC2148686F2B562665C3891507E35 (I288F847370AB993102C86AB98BD79E53 [0]),
.ICDAEEEBA9B4A4C5EBF042C0215A7BB0E (ID39228DB5F904D97CC6F69301B95F2D9 )); IEF91D04B90E6EC355FF6DD49C50BA7EA ICFAEEDAFB0F237713BE626AABCA45EE1 (.I7694F4A66316E53C8CDD9D9954BD611D (I288F847370AB993102C86AB98BD79E53 [2]),
.I0A3BC2148686F2B562665C3891507E35 (I288F847370AB993102C86AB98BD79E53 [1]), .ICDAEEEBA9B4A4C5EBF042C0215A7BB0E (ID39228DB5F904D97CC6F69301B95F2D9 )); IEF91D04B90E6EC355FF6DD49C50BA7EA
IF500A9C2C56DEBF8C12CA8C4E4895A29 (.I7694F4A66316E53C8CDD9D9954BD611D (I288F847370AB993102C86AB98BD79E53 [3]), .I0A3BC2148686F2B562665C3891507E35 (I288F847370AB993102C86AB98BD79E53 [2]),
.ICDAEEEBA9B4A4C5EBF042C0215A7BB0E (ID39228DB5F904D97CC6F69301B95F2D9 )); assign I975E762C6BF4B17F34E0966F54272008
= I76A88EC8C7A9140348BA5E2DAEEC0E89 ; wire I3B3DFD07FD7A0C6D0B4558504A4F6717 ; assign I3B3DFD07FD7A0C6D0B4558504A4F6717
= I8DE2A9CF71BCBDDB6996310B6090B645 ; reg [6:0] I02F288D1B97827548C2A777584D3E16E ; always @ (posedge I8DE2A9CF71BCBDDB6996310B6090B645 ) if (I975E762C6BF4B17F34E0966F54272008 ) I02F288D1B97827548C2A777584D3E16E
<= I37D350E5B2683ED4E78F696D8B080140 ; reg [3:0] IEF363218DA9C932A22163FA16CB46413 [6:0]; generate genvar I8CE4B16B22B58894AA86C421E8759DF3 ; for
(I8CE4B16B22B58894AA86C421E8759DF3 =0; I8CE4B16B22B58894AA86C421E8759DF3 <7; I8CE4B16B22B58894AA86C421E8759DF3 =I8CE4B16B22B58894AA86C421E8759DF3 +1) begin
: I41287185BB9B75BA2031272BB753FEBB wire ID674DFCD8B4DB6762BCB3667316D3BB9 , I9CFEFED8FB9497BAA5CD519D7D2BB5D7 ; assign
ID674DFCD8B4DB6762BCB3667316D3BB9 = I37D350E5B2683ED4E78F696D8B080140 [I8CE4B16B22B58894AA86C421E8759DF3 ] & ICFE6055D2E0503BE378BB63449EC7BA6 ;
assign I9CFEFED8FB9497BAA5CD519D7D2BB5D7 = I02F288D1B97827548C2A777584D3E16E [I8CE4B16B22B58894AA86C421E8759DF3 ]
& I0D28BD8A8650B66243673EBB8D515084 ; always @(posedge I3B3DFD07FD7A0C6D0B4558504A4F6717 ) begin if (I9CFEFED8FB9497BAA5CD519D7D2BB5D7 ) IEF363218DA9C932A22163FA16CB46413 [I8CE4B16B22B58894AA86C421E8759DF3 ]
<= I288F847370AB993102C86AB98BD79E53 ; else if (ID674DFCD8B4DB6762BCB3667316D3BB9 ) begin if (I76A88EC8C7A9140348BA5E2DAEEC0E89 ) IEF363218DA9C932A22163FA16CB46413 [I8CE4B16B22B58894AA86C421E8759DF3 ]
<= 4'd14; else IEF363218DA9C932A22163FA16CB46413 [I8CE4B16B22B58894AA86C421E8759DF3 ] <= 4'd15; end end end endgenerate
wire [3:0] IE458C04956F5B34B056E6C60536811A2 [6:0]; generate genvar I6F8F57715090DA2632453988D9A1501B ; for (I6F8F57715090DA2632453988D9A1501B =0;
I6F8F57715090DA2632453988D9A1501B <7; I6F8F57715090DA2632453988D9A1501B =I6F8F57715090DA2632453988D9A1501B +1) begin
: IF71B3896CAB4491397AAB7D180131EDA if ( I6F8F57715090DA2632453988D9A1501B ==0 ) assign IE458C04956F5B34B056E6C60536811A2 [I6F8F57715090DA2632453988D9A1501B ]
= IEF363218DA9C932A22163FA16CB46413 [I6F8F57715090DA2632453988D9A1501B ] & {4{IECAE13117D6F0584C25A9DA6C8F8415E [I6F8F57715090DA2632453988D9A1501B ]}}; else assign
IE458C04956F5B34B056E6C60536811A2 [I6F8F57715090DA2632453988D9A1501B ] = ( IEF363218DA9C932A22163FA16CB46413 [I6F8F57715090DA2632453988D9A1501B ]
& {4{IECAE13117D6F0584C25A9DA6C8F8415E [I6F8F57715090DA2632453988D9A1501B ]}} ) | IE458C04956F5B34B056E6C60536811A2 [I6F8F57715090DA2632453988D9A1501B -1]; end endgenerate
assign I8D777F385D3DFEC8815D20F7496026DC = IE458C04956F5B34B056E6C60536811A2 [6]; endmodule module IB51AA32163492596ADA06B22A9206E8F (I0A3BC2148686F2B562665C3891507E35 ,
I86266EE937D97F812A8E57D22B62EE29 , I27E9DD9482B253AA850544215471D9D5 , IE9DED2DF97E91174FD62E40E248B137D , I8715FEDE1A202C700CD025C90F3B2421 ,
I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 , IFC240E6D824E08568AA642A34947FEBC , I5844CE4E8F912137CD0A723AA7A4EBB2 , IF7F7CFDB9A31998C4AEFDC5C8BD5937A ,
IC68BD984558E67927B382A860837C32F , I47FE879774A01F989D46EFF34BCF4D44 , I1A7B4E094F07B0C85C5ACADEC807841F , I0F3FCCC5995F6CBAD0568AFF03FA9E41 ,
I082A499B7DDEF3C7897AB842B431A8AD , I89C5B8F33C91378743762C771A89F8C4 , I8357B924AEFCA0FDD29AADC1ABE078FF , I21345BCEA5A3A0213882E3493F7CE8A2 ,
IE8F9438C61FEFC48890126E846737803 , I00D170E901FDFA8C4D428ECAC839A4AB , I453DD3088EE862556BDD0F58B390F41F , I182E80B21C5A5F086FE70D9A01554365 ,
I346A81471C889B6C72A88423EB28B21A , I0EB8CC186C9B38B7FB99E477EE981265 , IF41F5F2D34464C2F1512CE4A38EAD286 , I75D612F1AEBBE1DC3FC1AC2ED5C21E7F ,
IA882574F5206B0DBAB0B61BA8B369A15 , IE78AFF6FF490ECAC5AFE4B8DF2BDC999 , I24D24CDA7F2D8B539E4F5C420BD826D9 , I61BAAAAF32AC5A7B6FFEBFC244A2D739 ,
I6E03B4F12533CBA29903F1C9DD1E5C3D , IAB9D6A507309488CCF13DB3F67F81B63 , I83FCEFDFE9F9D1C28AB321626447799F , I1905DD05FA116073F500B593198EED1C ,
I61E6EBA71A6BFA5A8FE92AB8FABECBBC , I79EB40C7CC07F0A913BA2E8F9D56D33B , I973092C325E8C2AE92FFF50B0288E777 , IB9445BEC437AE377554E2723C22C52B2 ,
I6A45CBE320E935B06BB0F08ECF1179D4 , I0EE48206D3023D05A5AA46FD33711C98 , I81414FA30C7BC73A9A778574097A714B , I4C39D6D4449338A7DA014742DE16FD46 ,
ID8E8746A568679217650DF444D98F91E , I30CD5687FB19DAD9CFD43FE994021B00 , I018477AF087A1484F83E54C386C2EF07 , I6970ADE3C1C5CEF4BF2ADF425B8B73CB ,
I4021D2C4A029457D9671036AF92F0AB8 , I6ABED3933223BDB35402C9F56973AB09 , I371CC04BDE216A35CEFED5553951955B , I032B17AEE0B7BC21B073F5A5AF886D30 ,
I64571D3B8AD6548BEF3F326B0C79154D , I528FBBEA2163A7F08F8CE87A6486A505 , IFD2E2FBE657226AA9EB0B69C70CEDAF0 , I6034EE230C5F2EA0D0828112861916C6 ,
I7E211F728072FEA639172DFD7FC475D2 , I4D5E955D6CD9D5E25ED4CE64CF4DC635 , I94F01074D91205FEBB9204892C80718F , IAE766072895E2EB8B8716944E133AE63 ); input
[0:1] IF7F7CFDB9A31998C4AEFDC5C8BD5937A , IC68BD984558E67927B382A860837C32F ; input wire I27E9DD9482B253AA850544215471D9D5 ,
I86266EE937D97F812A8E57D22B62EE29 ,I0A3BC2148686F2B562665C3891507E35 , I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 ; input
wire I47FE879774A01F989D46EFF34BCF4D44 ; output wire I1A7B4E094F07B0C85C5ACADEC807841F ; input [15:0] IFC240E6D824E08568AA642A34947FEBC ; output
[15:0] I5844CE4E8F912137CD0A723AA7A4EBB2 ; wire [15:0] I8D777F385D3DFEC8815D20F7496026DC ; input wire [3:0] IE9DED2DF97E91174FD62E40E248B137D ,
I8715FEDE1A202C700CD025C90F3B2421 ; input wire [8:0] I082A499B7DDEF3C7897AB842B431A8AD , I89C5B8F33C91378743762C771A89F8C4 ; input
wire [1:0] I8357B924AEFCA0FDD29AADC1ABE078FF ; input wire I21345BCEA5A3A0213882E3493F7CE8A2 , I00D170E901FDFA8C4D428ECAC839A4AB ,
IE8F9438C61FEFC48890126E846737803 ; input wire [1:0] I453DD3088EE862556BDD0F58B390F41F ; input wire [3:0] I182E80B21C5A5F086FE70D9A01554365 ; input
IF41F5F2D34464C2F1512CE4A38EAD286 , I75D612F1AEBBE1DC3FC1AC2ED5C21E7F , IA882574F5206B0DBAB0B61BA8B369A15 ; input
I346A81471C889B6C72A88423EB28B21A , I0EB8CC186C9B38B7FB99E477EE981265 ; output wire IE78AFF6FF490ECAC5AFE4B8DF2BDC999 ,
I24D24CDA7F2D8B539E4F5C420BD826D9 ; inout I61BAAAAF32AC5A7B6FFEBFC244A2D739 , I6E03B4F12533CBA29903F1C9DD1E5C3D ,
IAB9D6A507309488CCF13DB3F67F81B63 , I83FCEFDFE9F9D1C28AB321626447799F , I1905DD05FA116073F500B593198EED1C , I61E6EBA71A6BFA5A8FE92AB8FABECBBC ,
I79EB40C7CC07F0A913BA2E8F9D56D33B , I973092C325E8C2AE92FFF50B0288E777 , IB9445BEC437AE377554E2723C22C52B2 , I6A45CBE320E935B06BB0F08ECF1179D4 ,
I0EE48206D3023D05A5AA46FD33711C98 ; inout I81414FA30C7BC73A9A778574097A714B , I4C39D6D4449338A7DA014742DE16FD46 ,
ID8E8746A568679217650DF444D98F91E , I30CD5687FB19DAD9CFD43FE994021B00 , I018477AF087A1484F83E54C386C2EF07 , I6970ADE3C1C5CEF4BF2ADF425B8B73CB ,
I4021D2C4A029457D9671036AF92F0AB8 , I6ABED3933223BDB35402C9F56973AB09 , I371CC04BDE216A35CEFED5553951955B , I032B17AEE0B7BC21B073F5A5AF886D30 ,
I64571D3B8AD6548BEF3F326B0C79154D ; inout I528FBBEA2163A7F08F8CE87A6486A505 , IFD2E2FBE657226AA9EB0B69C70CEDAF0 ,
I6034EE230C5F2EA0D0828112861916C6 , I7E211F728072FEA639172DFD7FC475D2 , I4D5E955D6CD9D5E25ED4CE64CF4DC635 , I94F01074D91205FEBB9204892C80718F ; output
wire [1:0] IAE766072895E2EB8B8716944E133AE63 ; wire IAC0599EE2B1FB01124368C642A025AE6 , IB925B234F44A800CC3CE3166339BFB19 ; wire
[3:0] IB78E4CC26FAE6F795B778DAF30B00833 , ICDB60380CAC7C156C851A1AED5F82B18 ; assign IAC0599EE2B1FB01124368C642A025AE6
= I86266EE937D97F812A8E57D22B62EE29 ; assign IB925B234F44A800CC3CE3166339BFB19 = I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 ; assign
IB78E4CC26FAE6F795B778DAF30B00833 = IE9DED2DF97E91174FD62E40E248B137D ; assign ICDB60380CAC7C156C851A1AED5F82B18
= I8715FEDE1A202C700CD025C90F3B2421 ; wire [3:0] I975E762C6BF4B17F34E0966F54272008 ; wire [6:0] I37D350E5B2683ED4E78F696D8B080140 ;
wire [6:0] I2E16A98876DFFD2828D08E55F108424E ; wire ICFE6055D2E0503BE378BB63449EC7BA6 ; assign ICFE6055D2E0503BE378BB63449EC7BA6
= |I975E762C6BF4B17F34E0966F54272008 ; wire [3:0][3:0] I2E3034A0E1D9160A353BFB66B1405442 ; wire I6F2925832AC361C55FBABB66FC50F914 ; wire
[15:0] I51447734588298C46BA929BDC4DB0B94 ; assign I51447734588298C46BA929BDC4DB0B94 = {I2E3034A0E1D9160A353BFB66B1405442 [3],
I2E3034A0E1D9160A353BFB66B1405442 [2], I2E3034A0E1D9160A353BFB66B1405442 [1], I2E3034A0E1D9160A353BFB66B1405442 [0]}; wire
IC2E71DCCDB6779F28A7521AE60E49424 ; wire ID07E689D41DEE0A6E64AAFFE659AF67C ; assign IC2E71DCCDB6779F28A7521AE60E49424
= ID07E689D41DEE0A6E64AAFFE659AF67C & ~I6F2925832AC361C55FBABB66FC50F914 ; assign I8D777F385D3DFEC8815D20F7496026DC
= IC2E71DCCDB6779F28A7521AE60E49424 ? I51447734588298C46BA929BDC4DB0B94 : 0; assign I5844CE4E8F912137CD0A723AA7A4EBB2
= IFC240E6D824E08568AA642A34947FEBC | I8D777F385D3DFEC8815D20F7496026DC ; wire IB7F7EEB01501613F4B96A4710D3C8906 ; assign
IB7F7EEB01501613F4B96A4710D3C8906 = I0A3BC2148686F2B562665C3891507E35 & ~I6F2925832AC361C55FBABB66FC50F914 ; output
I0F3FCCC5995F6CBAD0568AFF03FA9E41 ; wire ID6299EFF2098B99E8BB408F652A2EE38 ; wire [0:1] IC9A7CC4AB393A8BD2AE6914033F0530B ,
ID78F9120B5CAEC4D064AF1B7C0EFA923 ; wire [0:1] I6EC93635F8FAC09674356349D7B864AB , I4B5D9EA056801D3FF5809343C7BC21C8 ; wire
[0:1] I882F749DD68DFEDCCCAC8ABDE84B58A5 , IDA4044D79AA1ECA013D47CA6A4D1D6B3 ; wire IAC00200163D6B8044E5259431846D3F8 ; wire
I149C2EAA6B8C9486634F6D592002E049 ; wire [3:0] IABF702906F6941BE8B9A1C1FAC6EED0F , IAAEEA8688711031D90BFAA8C7244F5E3 ; wire
IA387AEA270A27BDD008454099584DC16 , ICE66723AB312F38DC7058D59E9C120B4 ; I89B5FE0A834B8CEFBAD7FEA7A3D23364 IF5FA84218886B04F22503B6674ECC2D4 ( .IF41F5F2D34464C2F1512CE4A38EAD286 (IF41F5F2D34464C2F1512CE4A38EAD286 ),
.I75D612F1AEBBE1DC3FC1AC2ED5C21E7F (I75D612F1AEBBE1DC3FC1AC2ED5C21E7F ), .IA882574F5206B0DBAB0B61BA8B369A15 (IA882574F5206B0DBAB0B61BA8B369A15 ),
.I0EB8CC186C9B38B7FB99E477EE981265 (I0EB8CC186C9B38B7FB99E477EE981265 ), .IE78AFF6FF490ECAC5AFE4B8DF2BDC999 (IA387AEA270A27BDD008454099584DC16 ), .I21345BCEA5A3A0213882E3493F7CE8A2 (I21345BCEA5A3A0213882E3493F7CE8A2 ),
.IE8F9438C61FEFC48890126E846737803 (IE8F9438C61FEFC48890126E846737803 ), .I00D170E901FDFA8C4D428ECAC839A4AB (I00D170E901FDFA8C4D428ECAC839A4AB ), .I182E80B21C5A5F086FE70D9A01554365 (I182E80B21C5A5F086FE70D9A01554365 ),
.I453DD3088EE862556BDD0F58B390F41F (I453DD3088EE862556BDD0F58B390F41F ), .I346A81471C889B6C72A88423EB28B21A (I346A81471C889B6C72A88423EB28B21A ), .IABEB1D6F727D4016CBA8D230E06173E2 (I6EC93635F8FAC09674356349D7B864AB [0]), .IF365BCF55686BCCD839FE1624DD7D486 (IAC00200163D6B8044E5259431846D3F8 ),
.I5FBB67CECBAEE3FB61298BB458246F95 (I149C2EAA6B8C9486634F6D592002E049 ), .IDF6B1552FD717A0BD463ABC2AE6BE59A (IABF702906F6941BE8B9A1C1FAC6EED0F ),
.I10F9F36D10F50952745A860C2309B5EB (IAAEEA8688711031D90BFAA8C7244F5E3 ), .I9415662DEE73FC21C95CE7FCC2E8169E (IC9A7CC4AB393A8BD2AE6914033F0530B [0]),
.I24D24CDA7F2D8B539E4F5C420BD826D9 (ICE66723AB312F38DC7058D59E9C120B4 ) ); I55A61D3ABA6414EC766E337297B57941 IA31FCA8C33C497B87B9605EF487137F3 ( .I13B5BFE96F3E2FE411C9F66F4A582ADF (IF7F7CFDB9A31998C4AEFDC5C8BD5937A [0]),
.IEE02423CF012CD7FA6BC55B5769478E0 (I149C2EAA6B8C9486634F6D592002E049 ), .I55A302BB3928E3282F29EEAE2E18EC2F (I882F749DD68DFEDCCCAC8ABDE84B58A5 [0]),
.IF365BCF55686BCCD839FE1624DD7D486 (IAC00200163D6B8044E5259431846D3F8 ), .IDF6B1552FD717A0BD463ABC2AE6BE59A (IABF702906F6941BE8B9A1C1FAC6EED0F ),
.I10F9F36D10F50952745A860C2309B5EB (IAAEEA8688711031D90BFAA8C7244F5E3 ), .IF962DDDFCFB59F7648E592F6EAE19C93 (I61BAAAAF32AC5A7B6FFEBFC244A2D739 ),
.I0ED2ADDC6F83E144925F05986E9CFF86 (I6E03B4F12533CBA29903F1C9DD1E5C3D ), .IA95AE92E4828AF7B0DADD49D537FEE5E (IAB9D6A507309488CCF13DB3F67F81B63 ),
.I958F38294CE0C6337C616E28CE0C0EF4 (I83FCEFDFE9F9D1C28AB321626447799F ), .I531D5C1FBCF6E356CAFEEBA55A5B73D0 (I1905DD05FA116073F500B593198EED1C ),
.I3405A5272BCD250BE6AAB2071FA8E2C7 (I61E6EBA71A6BFA5A8FE92AB8FABECBBC ), .I0F71A3473EE22B4B3DACA05365112EB4 (I79EB40C7CC07F0A913BA2E8F9D56D33B ),
.IE3B0A4C4EA55DD2B44B6B72D7B0966A2 (I973092C325E8C2AE92FFF50B0288E777 ), .I2F93BC5D4AA9CC738D29F51E46D80581 (IB9445BEC437AE377554E2723C22C52B2 ),
.I6F8FB1BAF897A3508E8CE28CC0047AFE (I6A45CBE320E935B06BB0F08ECF1179D4 ), .I5E982716C925AA53DFAD54323E066CD2 (I0EE48206D3023D05A5AA46FD33711C98 ), .IEC862DB7074FDEA6C45E0A9D0E0686AA (I4D5E955D6CD9D5E25ED4CE64CF4DC635 ),
.I93C3BBEFFBA9F812B4F648566A44CBF6 (I6034EE230C5F2EA0D0828112861916C6 ), .I9BDAB36ABD4002A5BA799112841E27EE (I528FBBEA2163A7F08F8CE87A6486A505 ),
.ICB08DEE97A30C2949B48D36FB3C13CDC (), .IFAF919B89CA534E031F1812006C3375A (), .IDBE396CC46DEA10B12BE45753CAF92DD (),
.I074D81A9C803372CDEF5EF96C7A2E0BE (), .I441F445D5DBBC34DBE59585BE4CF0255 (), .IC056EF971E478FC69154775A88683389 (),
.I24FE5443C8249835AA81176E50160B25 () ); I6CCBE3F36B144174D7B5131F1612067F IBE369F38582F4AE93153D35BB7CE573C ( .IABEB1D6F727D4016CBA8D230E06173E2 (IC9A7CC4AB393A8BD2AE6914033F0530B [0]),
.I975E762C6BF4B17F34E0966F54272008 (I975E762C6BF4B17F34E0966F54272008 [0]), .I37D350E5B2683ED4E78F696D8B080140 (I37D350E5B2683ED4E78F696D8B080140 ), .ICFE6055D2E0503BE378BB63449EC7BA6 (ICFE6055D2E0503BE378BB63449EC7BA6 ), .IECAE13117D6F0584C25A9DA6C8F8415E (I2E16A98876DFFD2828D08E55F108424E ), .I8D777F385D3DFEC8815D20F7496026DC (I2E3034A0E1D9160A353BFB66B1405442 [0]), .I0A3BC2148686F2B562665C3891507E35 (IB7F7EEB01501613F4B96A4710D3C8906 ),
.I86266EE937D97F812A8E57D22B62EE29 (IAC0599EE2B1FB01124368C642A025AE6 ), .ID6299EFF2098B99E8BB408F652A2EE38 (!ID6299EFF2098B99E8BB408F652A2EE38 ), .I4CA8F5C40F80B904A3A115368EF165BF (), .I8357B924AEFCA0FDD29AADC1ABE078FF (I8357B924AEFCA0FDD29AADC1ABE078FF ) ); wire
I3882FD3F3EE3FD3421D92854F89E9B74 ; wire I056CD83F692E935A083F279DB3E4A49B ; wire [3:0] I46534ACB4986315DA02BC254874ABC07 ,
I282B6D08C46D42D08D98DE1F1981F108 ; wire ICFA37EB2734833DA0CD9A42455B20407 , I0B323720B6C803E4A14BFDB815005A25 ; I89B5FE0A834B8CEFBAD7FEA7A3D23364
I3E6741E20069866CF884E684771AC472 ( .IF41F5F2D34464C2F1512CE4A38EAD286 (IF41F5F2D34464C2F1512CE4A38EAD286 ), .I75D612F1AEBBE1DC3FC1AC2ED5C21E7F (I75D612F1AEBBE1DC3FC1AC2ED5C21E7F ),
.IA882574F5206B0DBAB0B61BA8B369A15 (IA387AEA270A27BDD008454099584DC16 ), .I0EB8CC186C9B38B7FB99E477EE981265 (I0EB8CC186C9B38B7FB99E477EE981265 ),
.IE78AFF6FF490ECAC5AFE4B8DF2BDC999 (ICFA37EB2734833DA0CD9A42455B20407 ), .I21345BCEA5A3A0213882E3493F7CE8A2 (I21345BCEA5A3A0213882E3493F7CE8A2 ),
.IE8F9438C61FEFC48890126E846737803 (IE8F9438C61FEFC48890126E846737803 ), .I00D170E901FDFA8C4D428ECAC839A4AB (I00D170E901FDFA8C4D428ECAC839A4AB ), .I182E80B21C5A5F086FE70D9A01554365 (I182E80B21C5A5F086FE70D9A01554365 ),
.I453DD3088EE862556BDD0F58B390F41F (I453DD3088EE862556BDD0F58B390F41F ), .I346A81471C889B6C72A88423EB28B21A (I346A81471C889B6C72A88423EB28B21A ), .IABEB1D6F727D4016CBA8D230E06173E2 (I6EC93635F8FAC09674356349D7B864AB [1]), .IF365BCF55686BCCD839FE1624DD7D486 (I3882FD3F3EE3FD3421D92854F89E9B74 ),
.I5FBB67CECBAEE3FB61298BB458246F95 (I056CD83F692E935A083F279DB3E4A49B ), .IDF6B1552FD717A0BD463ABC2AE6BE59A (I46534ACB4986315DA02BC254874ABC07 ),
.I10F9F36D10F50952745A860C2309B5EB (I282B6D08C46D42D08D98DE1F1981F108 ), .I9415662DEE73FC21C95CE7FCC2E8169E (IC9A7CC4AB393A8BD2AE6914033F0530B [1]),
.I24D24CDA7F2D8B539E4F5C420BD826D9 (I0B323720B6C803E4A14BFDB815005A25 ) ); I55A61D3ABA6414EC766E337297B57941 IF9F679C1B330AF90DA5CDA656066AD2D ( .I13B5BFE96F3E2FE411C9F66F4A582ADF (IF7F7CFDB9A31998C4AEFDC5C8BD5937A [1]),
.IEE02423CF012CD7FA6BC55B5769478E0 (I056CD83F692E935A083F279DB3E4A49B ), .I55A302BB3928E3282F29EEAE2E18EC2F (I882F749DD68DFEDCCCAC8ABDE84B58A5 [1]),
.IF365BCF55686BCCD839FE1624DD7D486 (I3882FD3F3EE3FD3421D92854F89E9B74 ), .IDF6B1552FD717A0BD463ABC2AE6BE59A (I46534ACB4986315DA02BC254874ABC07 ),
.I10F9F36D10F50952745A860C2309B5EB (I282B6D08C46D42D08D98DE1F1981F108 ), .IF962DDDFCFB59F7648E592F6EAE19C93 (I61BAAAAF32AC5A7B6FFEBFC244A2D739 ),
.I0ED2ADDC6F83E144925F05986E9CFF86 (I6E03B4F12533CBA29903F1C9DD1E5C3D ), .IA95AE92E4828AF7B0DADD49D537FEE5E (IAB9D6A507309488CCF13DB3F67F81B63 ),
.I958F38294CE0C6337C616E28CE0C0EF4 (I83FCEFDFE9F9D1C28AB321626447799F ), .I531D5C1FBCF6E356CAFEEBA55A5B73D0 (I1905DD05FA116073F500B593198EED1C ),
.I3405A5272BCD250BE6AAB2071FA8E2C7 (I61E6EBA71A6BFA5A8FE92AB8FABECBBC ), .I0F71A3473EE22B4B3DACA05365112EB4 (I79EB40C7CC07F0A913BA2E8F9D56D33B ),
.IE3B0A4C4EA55DD2B44B6B72D7B0966A2 (I973092C325E8C2AE92FFF50B0288E777 ), .I2F93BC5D4AA9CC738D29F51E46D80581 (IB9445BEC437AE377554E2723C22C52B2 ),
.I6F8FB1BAF897A3508E8CE28CC0047AFE (I6A45CBE320E935B06BB0F08ECF1179D4 ), .I5E982716C925AA53DFAD54323E066CD2 (I0EE48206D3023D05A5AA46FD33711C98 ), .IEC862DB7074FDEA6C45E0A9D0E0686AA (),
.I93C3BBEFFBA9F812B4F648566A44CBF6 (), .I9BDAB36ABD4002A5BA799112841E27EE (), .ICB08DEE97A30C2949B48D36FB3C13CDC (),
.IFAF919B89CA534E031F1812006C3375A (), .IDBE396CC46DEA10B12BE45753CAF92DD (), .I074D81A9C803372CDEF5EF96C7A2E0BE (),
.I441F445D5DBBC34DBE59585BE4CF0255 (), .IC056EF971E478FC69154775A88683389 (), .I24FE5443C8249835AA81176E50160B25 () ); I6CCBE3F36B144174D7B5131F1612067F
I2F39D4C17F5F2296550FBEDACEFB5C6C ( .IABEB1D6F727D4016CBA8D230E06173E2 (IC9A7CC4AB393A8BD2AE6914033F0530B [1]),
.I975E762C6BF4B17F34E0966F54272008 (I975E762C6BF4B17F34E0966F54272008 [1]), .I37D350E5B2683ED4E78F696D8B080140 (I37D350E5B2683ED4E78F696D8B080140 ), .ICFE6055D2E0503BE378BB63449EC7BA6 (ICFE6055D2E0503BE378BB63449EC7BA6 ), .IECAE13117D6F0584C25A9DA6C8F8415E (I2E16A98876DFFD2828D08E55F108424E ), .I8D777F385D3DFEC8815D20F7496026DC (I2E3034A0E1D9160A353BFB66B1405442 [1]), .I0A3BC2148686F2B562665C3891507E35 (IB7F7EEB01501613F4B96A4710D3C8906 ),
.I86266EE937D97F812A8E57D22B62EE29 (IAC0599EE2B1FB01124368C642A025AE6 ), .ID6299EFF2098B99E8BB408F652A2EE38 (!ID6299EFF2098B99E8BB408F652A2EE38 ), .I4CA8F5C40F80B904A3A115368EF165BF (), .I8357B924AEFCA0FDD29AADC1ABE078FF (I8357B924AEFCA0FDD29AADC1ABE078FF ) ); wire
I146DF6F0D72376116DDA3D656FCEDEF0 ; wire IE6BB1B855BD141D9BE228DF5B165F669 ; wire [3:0] I50879B1032EDCDD09F1DB7D9B88E6CF7 ,
I6C18BE9E78B5EF8AC5A74586B8515A12 ; wire I18FAF162006F440E660B7C2A52EDDA75 , I107EB23DABB0E9628572335AD5824055 ; I89B5FE0A834B8CEFBAD7FEA7A3D23364
I301FF87D9211990A754D0D3E0E8EFC08 ( .IF41F5F2D34464C2F1512CE4A38EAD286 (IF41F5F2D34464C2F1512CE4A38EAD286 ), .I75D612F1AEBBE1DC3FC1AC2ED5C21E7F (I75D612F1AEBBE1DC3FC1AC2ED5C21E7F ),
.IA882574F5206B0DBAB0B61BA8B369A15 (ICFA37EB2734833DA0CD9A42455B20407 ), .I0EB8CC186C9B38B7FB99E477EE981265 (I0EB8CC186C9B38B7FB99E477EE981265 ),
.IE78AFF6FF490ECAC5AFE4B8DF2BDC999 (I18FAF162006F440E660B7C2A52EDDA75 ), .I21345BCEA5A3A0213882E3493F7CE8A2 (I21345BCEA5A3A0213882E3493F7CE8A2 ),
.IE8F9438C61FEFC48890126E846737803 (IE8F9438C61FEFC48890126E846737803 ), .I00D170E901FDFA8C4D428ECAC839A4AB (I00D170E901FDFA8C4D428ECAC839A4AB ), .I182E80B21C5A5F086FE70D9A01554365 (I182E80B21C5A5F086FE70D9A01554365 ),
.I453DD3088EE862556BDD0F58B390F41F (I453DD3088EE862556BDD0F58B390F41F ), .I346A81471C889B6C72A88423EB28B21A (I346A81471C889B6C72A88423EB28B21A ), .IABEB1D6F727D4016CBA8D230E06173E2 (I4B5D9EA056801D3FF5809343C7BC21C8 [0]), .IF365BCF55686BCCD839FE1624DD7D486 (I146DF6F0D72376116DDA3D656FCEDEF0 ),
.I5FBB67CECBAEE3FB61298BB458246F95 (IE6BB1B855BD141D9BE228DF5B165F669 ), .IDF6B1552FD717A0BD463ABC2AE6BE59A (I50879B1032EDCDD09F1DB7D9B88E6CF7 ),
.I10F9F36D10F50952745A860C2309B5EB (I6C18BE9E78B5EF8AC5A74586B8515A12 ), .I9415662DEE73FC21C95CE7FCC2E8169E (ID78F9120B5CAEC4D064AF1B7C0EFA923 [0]),
.I24D24CDA7F2D8B539E4F5C420BD826D9 (I107EB23DABB0E9628572335AD5824055 ) ); I55A61D3ABA6414EC766E337297B57941 I85138BA82CA09CC9D0E7536D68EE9D08 ( .I13B5BFE96F3E2FE411C9F66F4A582ADF (IC68BD984558E67927B382A860837C32F [0]),
.IEE02423CF012CD7FA6BC55B5769478E0 (IE6BB1B855BD141D9BE228DF5B165F669 ), .I55A302BB3928E3282F29EEAE2E18EC2F (IDA4044D79AA1ECA013D47CA6A4D1D6B3 [0]),
.IF365BCF55686BCCD839FE1624DD7D486 (I146DF6F0D72376116DDA3D656FCEDEF0 ), .IDF6B1552FD717A0BD463ABC2AE6BE59A (I50879B1032EDCDD09F1DB7D9B88E6CF7 ),
.I10F9F36D10F50952745A860C2309B5EB (I6C18BE9E78B5EF8AC5A74586B8515A12 ), .IF962DDDFCFB59F7648E592F6EAE19C93 (I81414FA30C7BC73A9A778574097A714B ),
.I0ED2ADDC6F83E144925F05986E9CFF86 (I4C39D6D4449338A7DA014742DE16FD46 ), .IA95AE92E4828AF7B0DADD49D537FEE5E (ID8E8746A568679217650DF444D98F91E ),
.I958F38294CE0C6337C616E28CE0C0EF4 (I30CD5687FB19DAD9CFD43FE994021B00 ), .I531D5C1FBCF6E356CAFEEBA55A5B73D0 (I018477AF087A1484F83E54C386C2EF07 ),
.I3405A5272BCD250BE6AAB2071FA8E2C7 (I6970ADE3C1C5CEF4BF2ADF425B8B73CB ), .I0F71A3473EE22B4B3DACA05365112EB4 (I4021D2C4A029457D9671036AF92F0AB8 ),
.IE3B0A4C4EA55DD2B44B6B72D7B0966A2 (I6ABED3933223BDB35402C9F56973AB09 ), .I2F93BC5D4AA9CC738D29F51E46D80581 (I371CC04BDE216A35CEFED5553951955B ),
.I6F8FB1BAF897A3508E8CE28CC0047AFE (I032B17AEE0B7BC21B073F5A5AF886D30 ), .I5E982716C925AA53DFAD54323E066CD2 (I64571D3B8AD6548BEF3F326B0C79154D ), .IEC862DB7074FDEA6C45E0A9D0E0686AA (I94F01074D91205FEBB9204892C80718F ),
.I93C3BBEFFBA9F812B4F648566A44CBF6 (I7E211F728072FEA639172DFD7FC475D2 ), .I9BDAB36ABD4002A5BA799112841E27EE (IFD2E2FBE657226AA9EB0B69C70CEDAF0 ),
.ICB08DEE97A30C2949B48D36FB3C13CDC (), .IFAF919B89CA534E031F1812006C3375A (), .IDBE396CC46DEA10B12BE45753CAF92DD (),
.I074D81A9C803372CDEF5EF96C7A2E0BE (), .I441F445D5DBBC34DBE59585BE4CF0255 (), .IC056EF971E478FC69154775A88683389 (),
.I24FE5443C8249835AA81176E50160B25 () ); I6CCBE3F36B144174D7B5131F1612067F ID465F65225F0C42CEEF7697329CF83DD ( .IABEB1D6F727D4016CBA8D230E06173E2 (ID78F9120B5CAEC4D064AF1B7C0EFA923 [0]),
.I975E762C6BF4B17F34E0966F54272008 (I975E762C6BF4B17F34E0966F54272008 [2]), .I37D350E5B2683ED4E78F696D8B080140 (I37D350E5B2683ED4E78F696D8B080140 ), .ICFE6055D2E0503BE378BB63449EC7BA6 (ICFE6055D2E0503BE378BB63449EC7BA6 ), .IECAE13117D6F0584C25A9DA6C8F8415E (I2E16A98876DFFD2828D08E55F108424E ), .I8D777F385D3DFEC8815D20F7496026DC (I2E3034A0E1D9160A353BFB66B1405442 [2]), .I0A3BC2148686F2B562665C3891507E35 (IB7F7EEB01501613F4B96A4710D3C8906 ),
.I86266EE937D97F812A8E57D22B62EE29 (IAC0599EE2B1FB01124368C642A025AE6 ), .ID6299EFF2098B99E8BB408F652A2EE38 (!ID6299EFF2098B99E8BB408F652A2EE38 ), .I4CA8F5C40F80B904A3A115368EF165BF (), .I8357B924AEFCA0FDD29AADC1ABE078FF (I8357B924AEFCA0FDD29AADC1ABE078FF ) ); wire
I5C12871940B6DDB931295F6AB41E27A9 ; wire ID33ED9DAD0D654ECA586ACD097C0ECFC ; wire [3:0] I1341B411C8C289AABF48A9A2DCB1A23B ,
IDEE66ED5577CB6B7691E39CAB404366C ; wire IA45557FF6F2E75FCAD293F1A990F410E ; I89B5FE0A834B8CEFBAD7FEA7A3D23364 I44C8D082C06FF81F0EB37A2D6F1D4218 ( .IF41F5F2D34464C2F1512CE4A38EAD286 (IF41F5F2D34464C2F1512CE4A38EAD286 ),
.I75D612F1AEBBE1DC3FC1AC2ED5C21E7F (I75D612F1AEBBE1DC3FC1AC2ED5C21E7F ), .IA882574F5206B0DBAB0B61BA8B369A15 (I18FAF162006F440E660B7C2A52EDDA75 ),
.I0EB8CC186C9B38B7FB99E477EE981265 (I0EB8CC186C9B38B7FB99E477EE981265 ), .IE78AFF6FF490ECAC5AFE4B8DF2BDC999 (IE78AFF6FF490ECAC5AFE4B8DF2BDC999 ), .I21345BCEA5A3A0213882E3493F7CE8A2 (I21345BCEA5A3A0213882E3493F7CE8A2 ),
.IE8F9438C61FEFC48890126E846737803 (IE8F9438C61FEFC48890126E846737803 ), .I00D170E901FDFA8C4D428ECAC839A4AB (I00D170E901FDFA8C4D428ECAC839A4AB ), .I182E80B21C5A5F086FE70D9A01554365 (I182E80B21C5A5F086FE70D9A01554365 ),
.I453DD3088EE862556BDD0F58B390F41F (I453DD3088EE862556BDD0F58B390F41F ), .I346A81471C889B6C72A88423EB28B21A (I346A81471C889B6C72A88423EB28B21A ), .IABEB1D6F727D4016CBA8D230E06173E2 (I4B5D9EA056801D3FF5809343C7BC21C8 [1]), .IF365BCF55686BCCD839FE1624DD7D486 (I5C12871940B6DDB931295F6AB41E27A9 ),
.I5FBB67CECBAEE3FB61298BB458246F95 (ID33ED9DAD0D654ECA586ACD097C0ECFC ), .IDF6B1552FD717A0BD463ABC2AE6BE59A (I1341B411C8C289AABF48A9A2DCB1A23B ),
.I10F9F36D10F50952745A860C2309B5EB (IDEE66ED5577CB6B7691E39CAB404366C ), .I9415662DEE73FC21C95CE7FCC2E8169E (ID78F9120B5CAEC4D064AF1B7C0EFA923 [1]),
.I24D24CDA7F2D8B539E4F5C420BD826D9 (IA45557FF6F2E75FCAD293F1A990F410E ) ); I55A61D3ABA6414EC766E337297B57941 I45D78A8C0A32B9DC806FC6446F5F7FA8 ( .I13B5BFE96F3E2FE411C9F66F4A582ADF (IC68BD984558E67927B382A860837C32F [1]),
.IEE02423CF012CD7FA6BC55B5769478E0 (ID33ED9DAD0D654ECA586ACD097C0ECFC ), .I55A302BB3928E3282F29EEAE2E18EC2F (IDA4044D79AA1ECA013D47CA6A4D1D6B3 [1]),
.IF365BCF55686BCCD839FE1624DD7D486 (I5C12871940B6DDB931295F6AB41E27A9 ), .IDF6B1552FD717A0BD463ABC2AE6BE59A (I1341B411C8C289AABF48A9A2DCB1A23B ),
.I10F9F36D10F50952745A860C2309B5EB (IDEE66ED5577CB6B7691E39CAB404366C ), .IF962DDDFCFB59F7648E592F6EAE19C93 (I81414FA30C7BC73A9A778574097A714B ),
.I0ED2ADDC6F83E144925F05986E9CFF86 (I4C39D6D4449338A7DA014742DE16FD46 ), .IA95AE92E4828AF7B0DADD49D537FEE5E (ID8E8746A568679217650DF444D98F91E ),
.I958F38294CE0C6337C616E28CE0C0EF4 (I30CD5687FB19DAD9CFD43FE994021B00 ), .I531D5C1FBCF6E356CAFEEBA55A5B73D0 (I018477AF087A1484F83E54C386C2EF07 ),
.I3405A5272BCD250BE6AAB2071FA8E2C7 (I6970ADE3C1C5CEF4BF2ADF425B8B73CB ), .I0F71A3473EE22B4B3DACA05365112EB4 (I4021D2C4A029457D9671036AF92F0AB8 ),
.IE3B0A4C4EA55DD2B44B6B72D7B0966A2 (I6ABED3933223BDB35402C9F56973AB09 ), .I2F93BC5D4AA9CC738D29F51E46D80581 (I371CC04BDE216A35CEFED5553951955B ),
.I6F8FB1BAF897A3508E8CE28CC0047AFE (I032B17AEE0B7BC21B073F5A5AF886D30 ), .I5E982716C925AA53DFAD54323E066CD2 (I64571D3B8AD6548BEF3F326B0C79154D ), .IEC862DB7074FDEA6C45E0A9D0E0686AA (),
.I93C3BBEFFBA9F812B4F648566A44CBF6 (), .I9BDAB36ABD4002A5BA799112841E27EE (), .ICB08DEE97A30C2949B48D36FB3C13CDC (),
.IFAF919B89CA534E031F1812006C3375A (), .IDBE396CC46DEA10B12BE45753CAF92DD (), .I074D81A9C803372CDEF5EF96C7A2E0BE (),
.I441F445D5DBBC34DBE59585BE4CF0255 (), .IC056EF971E478FC69154775A88683389 (), .I24FE5443C8249835AA81176E50160B25 () ); I6CCBE3F36B144174D7B5131F1612067F
I183C5AB93B7C78DB5E7CD0BD5591C481 ( .IABEB1D6F727D4016CBA8D230E06173E2 (ID78F9120B5CAEC4D064AF1B7C0EFA923 [1]),
.I975E762C6BF4B17F34E0966F54272008 (I975E762C6BF4B17F34E0966F54272008 [3]), .I37D350E5B2683ED4E78F696D8B080140 (I37D350E5B2683ED4E78F696D8B080140 ), .ICFE6055D2E0503BE378BB63449EC7BA6 (ICFE6055D2E0503BE378BB63449EC7BA6 ), .IECAE13117D6F0584C25A9DA6C8F8415E (I2E16A98876DFFD2828D08E55F108424E ), .I8D777F385D3DFEC8815D20F7496026DC (I2E3034A0E1D9160A353BFB66B1405442 [3]), .I0A3BC2148686F2B562665C3891507E35 (IB7F7EEB01501613F4B96A4710D3C8906 ),
.I86266EE937D97F812A8E57D22B62EE29 (IAC0599EE2B1FB01124368C642A025AE6 ), .ID6299EFF2098B99E8BB408F652A2EE38 (!ID6299EFF2098B99E8BB408F652A2EE38 ), .I4CA8F5C40F80B904A3A115368EF165BF (), .I8357B924AEFCA0FDD29AADC1ABE078FF (I8357B924AEFCA0FDD29AADC1ABE078FF ) ); I3A7EEC60129C000F5EF89FDB38307204
I6027381B66C3039F503013E521C6285B ( .ICFE6055D2E0503BE378BB63449EC7BA6 (ICFE6055D2E0503BE378BB63449EC7BA6 ), .I9EC4C0AFD450CEAC7ADB81C3BCFC9732 (I27E9DD9482B253AA850544215471D9D5 ),
.I86266EE937D97F812A8E57D22B62EE29 (IAC0599EE2B1FB01124368C642A025AE6 ), .I0A3BC2148686F2B562665C3891507E35 (IB7F7EEB01501613F4B96A4710D3C8906 ),
.I47FE879774A01F989D46EFF34BCF4D44 (I47FE879774A01F989D46EFF34BCF4D44 ), .I1A7B4E094F07B0C85C5ACADEC807841F (I1A7B4E094F07B0C85C5ACADEC807841F ),
.IB4CDA117A366592F9BB0BF24B8090648 (IB925B234F44A800CC3CE3166339BFB19 ), .I662D272D5B777249F5AD3F0BD29F079C (IB78E4CC26FAE6F795B778DAF30B00833 ), .I1653E44E546EA269CD4BEFADAFD0F53C (ICDB60380CAC7C156C851A1AED5F82B18 ), .IC28D2F5880CB3E1E4D819DD6223D52D5 (ID07E689D41DEE0A6E64AAFFE659AF67C ), .I37D350E5B2683ED4E78F696D8B080140 (I37D350E5B2683ED4E78F696D8B080140 ), .IECAE13117D6F0584C25A9DA6C8F8415E (I2E16A98876DFFD2828D08E55F108424E ), .I5EBEE840AC1BD9B012986A05E8BD96CC (I0F3FCCC5995F6CBAD0568AFF03FA9E41 ), .I5D66DC68084DBC91ECB34E334C1BC291 (I082A499B7DDEF3C7897AB842B431A8AD ), .I51E96C20C528EDDF5025F8B0F8448C53 (I89C5B8F33C91378743762C771A89F8C4 ), .I6F2925832AC361C55FBABB66FC50F914 (I6F2925832AC361C55FBABB66FC50F914 ) ); assign
I6F2925832AC361C55FBABB66FC50F914 = IAC00200163D6B8044E5259431846D3F8 & I3882FD3F3EE3FD3421D92854F89E9B74 & I146DF6F0D72376116DDA3D656FCEDEF0
& I5C12871940B6DDB931295F6AB41E27A9 ; assign I24D24CDA7F2D8B539E4F5C420BD826D9 = ICE66723AB312F38DC7058D59E9C120B4
| I0B323720B6C803E4A14BFDB815005A25 | I107EB23DABB0E9628572335AD5824055 | IA45557FF6F2E75FCAD293F1A990F410E ; assign
I4B5D9EA056801D3FF5809343C7BC21C8 = IDA4044D79AA1ECA013D47CA6A4D1D6B3 ; assign I6EC93635F8FAC09674356349D7B864AB
= I882F749DD68DFEDCCCAC8ABDE84B58A5 ; assign IAE766072895E2EB8B8716944E133AE63 [0] = !I4B5D9EA056801D3FF5809343C7BC21C8 [1]; assign
IAE766072895E2EB8B8716944E133AE63 [1] = !I4B5D9EA056801D3FF5809343C7BC21C8 [0]; endmodule module I55A61D3ABA6414EC766E337297B57941 (
input wire IF365BCF55686BCCD839FE1624DD7D486 , IEE02423CF012CD7FA6BC55B5769478E0 , input wire [3:0] IDF6B1552FD717A0BD463ABC2AE6BE59A ,
I10F9F36D10F50952745A860C2309B5EB , output wire I55A302BB3928E3282F29EEAE2E18EC2F , input wire I13B5BFE96F3E2FE411C9F66F4A582ADF , inout
wire IF962DDDFCFB59F7648E592F6EAE19C93 , I0ED2ADDC6F83E144925F05986E9CFF86 , IA95AE92E4828AF7B0DADD49D537FEE5E ,
I958F38294CE0C6337C616E28CE0C0EF4 , I531D5C1FBCF6E356CAFEEBA55A5B73D0 , I3405A5272BCD250BE6AAB2071FA8E2C7 , I0F71A3473EE22B4B3DACA05365112EB4 ,
IE3B0A4C4EA55DD2B44B6B72D7B0966A2 , I2F93BC5D4AA9CC738D29F51E46D80581 , I6F8FB1BAF897A3508E8CE28CC0047AFE , I5E982716C925AA53DFAD54323E066CD2 , inout
wire IEC862DB7074FDEA6C45E0A9D0E0686AA , inout wire I93C3BBEFFBA9F812B4F648566A44CBF6 , inout wire I9BDAB36ABD4002A5BA799112841E27EE , inout
wire ICB08DEE97A30C2949B48D36FB3C13CDC , inout wire IFAF919B89CA534E031F1812006C3375A , inout wire IDBE396CC46DEA10B12BE45753CAF92DD , inout
wire I074D81A9C803372CDEF5EF96C7A2E0BE , inout wire I441F445D5DBBC34DBE59585BE4CF0255 , inout wire IC056EF971E478FC69154775A88683389 , inout
wire I24FE5443C8249835AA81176E50160B25 ); wire I8FC22CBFEC954567F81E436DBF1AE83A ; assign I8FC22CBFEC954567F81E436DBF1AE83A
= I0ED2ADDC6F83E144925F05986E9CFF86 | IA95AE92E4828AF7B0DADD49D537FEE5E | I958F38294CE0C6337C616E28CE0C0EF4 | I531D5C1FBCF6E356CAFEEBA55A5B73D0
| I3405A5272BCD250BE6AAB2071FA8E2C7 | I0F71A3473EE22B4B3DACA05365112EB4 | IE3B0A4C4EA55DD2B44B6B72D7B0966A2 | I2F93BC5D4AA9CC738D29F51E46D80581
| I6F8FB1BAF897A3508E8CE28CC0047AFE | I5E982716C925AA53DFAD54323E066CD2 ; reg I86F2E62365A4DAB2D24CA8D4F6C1FBD3 ; assign
I55A302BB3928E3282F29EEAE2E18EC2F = ~( (I13B5BFE96F3E2FE411C9F66F4A582ADF | I86F2E62365A4DAB2D24CA8D4F6C1FBD3 )
& !IF365BCF55686BCCD839FE1624DD7D486 ) ;  initial begin I86F2E62365A4DAB2D24CA8D4F6C1FBD3 = 0; forever begin @(negedge
IF962DDDFCFB59F7648E592F6EAE19C93 ) I86F2E62365A4DAB2D24CA8D4F6C1FBD3 = I8FC22CBFEC954567F81E436DBF1AE83A & IEE02423CF012CD7FA6BC55B5769478E0 ; #(25*IDF6B1552FD717A0BD463ABC2AE6BE59A )
I86F2E62365A4DAB2D24CA8D4F6C1FBD3 = 0; end end endmodule module I379BDABA1FBE95FD8A49051997E9665F (I6F13D2E1112161FE6F8EA1EDD3F01310 ,
I208F156D4A803025C284BB595A7576B4 , I3F3B6F139F935CDE0338584380A06130 ); input wire I6F13D2E1112161FE6F8EA1EDD3F01310 ,
I208F156D4A803025C284BB595A7576B4 ; output wire I3F3B6F139F935CDE0338584380A06130 ; wire I9E8E4A3A68C2F178BE5AAAF290798A42 ; reg
IAEA5AEDB5A24E4DB6C6FC3D2FEA1E044 ; assign I9E8E4A3A68C2F178BE5AAAF290798A42 = ~I6F13D2E1112161FE6F8EA1EDD3F01310 ; always
@ (I9E8E4A3A68C2F178BE5AAAF290798A42 or I208F156D4A803025C284BB595A7576B4 ) if (I9E8E4A3A68C2F178BE5AAAF290798A42 ) IAEA5AEDB5A24E4DB6C6FC3D2FEA1E044
= I208F156D4A803025C284BB595A7576B4 ; assign I3F3B6F139F935CDE0338584380A06130 = I6F13D2E1112161FE6F8EA1EDD3F01310
& IAEA5AEDB5A24E4DB6C6FC3D2FEA1E044 ; endmodule module I9E18496CBD21D6A02574C0F31F3D3FB7 (I6F13D2E1112161FE6F8EA1EDD3F01310 ,
I208F156D4A803025C284BB595A7576B4 , I3F3B6F139F935CDE0338584380A06130 ); input wire I6F13D2E1112161FE6F8EA1EDD3F01310 ,I208F156D4A803025C284BB595A7576B4 ; output
wire I3F3B6F139F935CDE0338584380A06130 ; reg IAEA5AEDB5A24E4DB6C6FC3D2FEA1E044 ; always @ (I6F13D2E1112161FE6F8EA1EDD3F01310
or I208F156D4A803025C284BB595A7576B4 ) if (I6F13D2E1112161FE6F8EA1EDD3F01310 ) IAEA5AEDB5A24E4DB6C6FC3D2FEA1E044
= I208F156D4A803025C284BB595A7576B4 ; assign I3F3B6F139F935CDE0338584380A06130 = I6F13D2E1112161FE6F8EA1EDD3F01310
| ~IAEA5AEDB5A24E4DB6C6FC3D2FEA1E044 ; endmodule module I21F5A4F10878160CE707AC6682B91D1B (I2536792601E6CADEAB49502F1BD19044 , I27E9DD9482B253AA850544215471D9D5 ,
I86266EE937D97F812A8E57D22B62EE29 ,I0A3BC2148686F2B562665C3891507E35 , I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 , IE9DED2DF97E91174FD62E40E248B137D ,
I8715FEDE1A202C700CD025C90F3B2421 , I1A7B4E094F07B0C85C5ACADEC807841F , I21345BCEA5A3A0213882E3493F7CE8A2 , IE8F9438C61FEFC48890126E846737803 ,
I00D170E901FDFA8C4D428ECAC839A4AB , I453DD3088EE862556BDD0F58B390F41F , I182E80B21C5A5F086FE70D9A01554365 , I346A81471C889B6C72A88423EB28B21A ,
I0EB8CC186C9B38B7FB99E477EE981265 , IF41F5F2D34464C2F1512CE4A38EAD286 , I75D612F1AEBBE1DC3FC1AC2ED5C21E7F , IA882574F5206B0DBAB0B61BA8B369A15 ,
IE78AFF6FF490ECAC5AFE4B8DF2BDC999 , I24D24CDA7F2D8B539E4F5C420BD826D9 , I082A499B7DDEF3C7897AB842B431A8AD , I89C5B8F33C91378743762C771A89F8C4 ,
I8357B924AEFCA0FDD29AADC1ABE078FF , IF6068DAA29DBB05A7EAD1E3B5A48BBEE , IA70367AA7CB74E510F4F9413CCF059D3 , I61BAAAAF32AC5A7B6FFEBFC244A2D739 ,
I6E03B4F12533CBA29903F1C9DD1E5C3D , IAB9D6A507309488CCF13DB3F67F81B63 , I83FCEFDFE9F9D1C28AB321626447799F , I1905DD05FA116073F500B593198EED1C ,
I61E6EBA71A6BFA5A8FE92AB8FABECBBC , I79EB40C7CC07F0A913BA2E8F9D56D33B , I973092C325E8C2AE92FFF50B0288E777 , IB9445BEC437AE377554E2723C22C52B2 ,
I6A45CBE320E935B06BB0F08ECF1179D4 , I0EE48206D3023D05A5AA46FD33711C98 , I81414FA30C7BC73A9A778574097A714B , I4C39D6D4449338A7DA014742DE16FD46 ,
ID8E8746A568679217650DF444D98F91E , I30CD5687FB19DAD9CFD43FE994021B00 , I018477AF087A1484F83E54C386C2EF07 , I6970ADE3C1C5CEF4BF2ADF425B8B73CB ,
I4021D2C4A029457D9671036AF92F0AB8 , I6ABED3933223BDB35402C9F56973AB09 , I371CC04BDE216A35CEFED5553951955B , I032B17AEE0B7BC21B073F5A5AF886D30 ,
I64571D3B8AD6548BEF3F326B0C79154D , I5B9F987DBE3EDAC4E347A14A5782131F , I08C038534302D663980480E37D20BC83 , I769454D2A8D191F3E322B7B5DF928B5D ,
I01BDC194686F6DC3F502CFA733822312 , I87B3D78A5F6FFC46951ED28E772E594D , I159859469876028CEA112C7C16B1CAF5 , IAE766072895E2EB8B8716944E133AE63 ); localparam
I20215169A99BAB8B27571CCDC8331264 = 64; input wire [I20215169A99BAB8B27571CCDC8331264 *4-1:0] I2536792601E6CADEAB49502F1BD19044 ; input
wire I27E9DD9482B253AA850544215471D9D5 , I86266EE937D97F812A8E57D22B62EE29 ,I0A3BC2148686F2B562665C3891507E35 ,
I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 ; input wire [3:0] IE9DED2DF97E91174FD62E40E248B137D , I8715FEDE1A202C700CD025C90F3B2421 ; output
wire I1A7B4E094F07B0C85C5ACADEC807841F ; input wire [8:0] I082A499B7DDEF3C7897AB842B431A8AD , I89C5B8F33C91378743762C771A89F8C4 ; input
wire [1:0] I8357B924AEFCA0FDD29AADC1ABE078FF ; output wire [15:0] IF6068DAA29DBB05A7EAD1E3B5A48BBEE ; output wire
[5:0] IA70367AA7CB74E510F4F9413CCF059D3 ; input wire I21345BCEA5A3A0213882E3493F7CE8A2 , I00D170E901FDFA8C4D428ECAC839A4AB ,
IE8F9438C61FEFC48890126E846737803 ; input wire [1:0] I453DD3088EE862556BDD0F58B390F41F ; input wire [3:0] I182E80B21C5A5F086FE70D9A01554365 ; input
I346A81471C889B6C72A88423EB28B21A , I0EB8CC186C9B38B7FB99E477EE981265 ; input wire IF41F5F2D34464C2F1512CE4A38EAD286 ,
I75D612F1AEBBE1DC3FC1AC2ED5C21E7F , IA882574F5206B0DBAB0B61BA8B369A15 ; output wire IE78AFF6FF490ECAC5AFE4B8DF2BDC999 ,
I24D24CDA7F2D8B539E4F5C420BD826D9 ; inout wire [0:1] I61BAAAAF32AC5A7B6FFEBFC244A2D739 , I6E03B4F12533CBA29903F1C9DD1E5C3D ,
IAB9D6A507309488CCF13DB3F67F81B63 , I83FCEFDFE9F9D1C28AB321626447799F , I1905DD05FA116073F500B593198EED1C , I61E6EBA71A6BFA5A8FE92AB8FABECBBC ,
I79EB40C7CC07F0A913BA2E8F9D56D33B , I973092C325E8C2AE92FFF50B0288E777 , IB9445BEC437AE377554E2723C22C52B2 , I6A45CBE320E935B06BB0F08ECF1179D4 ,
I0EE48206D3023D05A5AA46FD33711C98 ; inout wire [0:1] I81414FA30C7BC73A9A778574097A714B , I4C39D6D4449338A7DA014742DE16FD46 ,
ID8E8746A568679217650DF444D98F91E , I30CD5687FB19DAD9CFD43FE994021B00 , I018477AF087A1484F83E54C386C2EF07 , I6970ADE3C1C5CEF4BF2ADF425B8B73CB ,
I4021D2C4A029457D9671036AF92F0AB8 , I6ABED3933223BDB35402C9F56973AB09 , I371CC04BDE216A35CEFED5553951955B , I032B17AEE0B7BC21B073F5A5AF886D30 ,
I64571D3B8AD6548BEF3F326B0C79154D ; inout wire [1:0] I5B9F987DBE3EDAC4E347A14A5782131F , I08C038534302D663980480E37D20BC83 ,
I769454D2A8D191F3E322B7B5DF928B5D , I01BDC194686F6DC3F502CFA733822312 , I87B3D78A5F6FFC46951ED28E772E594D , I159859469876028CEA112C7C16B1CAF5 ; output
wire [63:0] IAE766072895E2EB8B8716944E133AE63 ; wire [I20215169A99BAB8B27571CCDC8331264 *2-1:0] IC9A7CC4AB393A8BD2AE6914033F0530B ,
ID78F9120B5CAEC4D064AF1B7C0EFA923 ; assign IC9A7CC4AB393A8BD2AE6914033F0530B [I20215169A99BAB8B27571CCDC8331264 *2-1:I20215169A99BAB8B27571CCDC8331264 ]
= I2536792601E6CADEAB49502F1BD19044 [I20215169A99BAB8B27571CCDC8331264 *4-1:I20215169A99BAB8B27571CCDC8331264 *3]; assign
IC9A7CC4AB393A8BD2AE6914033F0530B [I20215169A99BAB8B27571CCDC8331264 -1:0] = I2536792601E6CADEAB49502F1BD19044 [I20215169A99BAB8B27571CCDC8331264 *2-1:I20215169A99BAB8B27571CCDC8331264 *1];
assign ID78F9120B5CAEC4D064AF1B7C0EFA923 [I20215169A99BAB8B27571CCDC8331264 *2-1:I20215169A99BAB8B27571CCDC8331264 ]
= I2536792601E6CADEAB49502F1BD19044 [I20215169A99BAB8B27571CCDC8331264 *3-1:I20215169A99BAB8B27571CCDC8331264 *2]; assign
ID78F9120B5CAEC4D064AF1B7C0EFA923 [I20215169A99BAB8B27571CCDC8331264 -1:0] = I2536792601E6CADEAB49502F1BD19044 [I20215169A99BAB8B27571CCDC8331264 *1-1:I20215169A99BAB8B27571CCDC8331264 *0]; wire
[15:0] ICE7D06150E11255C4F8EE2384429A32A [I20215169A99BAB8B27571CCDC8331264 :0]; assign ICE7D06150E11255C4F8EE2384429A32A [0]
= 0; assign IF6068DAA29DBB05A7EAD1E3B5A48BBEE = ICE7D06150E11255C4F8EE2384429A32A [I20215169A99BAB8B27571CCDC8331264 ]; wire
[I20215169A99BAB8B27571CCDC8331264 :0] IF8DEC8403A8BD60501F344A464CBF9AC ; assign IF8DEC8403A8BD60501F344A464CBF9AC [0]
= 0; assign I1A7B4E094F07B0C85C5ACADEC807841F = IF8DEC8403A8BD60501F344A464CBF9AC [I20215169A99BAB8B27571CCDC8331264 ]; wire
[I20215169A99BAB8B27571CCDC8331264 :0] IE22428CCF96CDA9674A939C209AD1000 ; assign IE22428CCF96CDA9674A939C209AD1000 [0]
= IA882574F5206B0DBAB0B61BA8B369A15 ; assign IE78AFF6FF490ECAC5AFE4B8DF2BDC999 = IE22428CCF96CDA9674A939C209AD1000 [I20215169A99BAB8B27571CCDC8331264 ]; wire
[I20215169A99BAB8B27571CCDC8331264 -1:0] I48A355561F0628CB2813BD54EADAA46C ; assign I24D24CDA7F2D8B539E4F5C420BD826D9
= |I48A355561F0628CB2813BD54EADAA46C ; reg I48F5E59356CCB45A1C41CAE764DF169C ; always @(I1A7B4E094F07B0C85C5ACADEC807841F
or I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 ) if ( I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 == 1'b0 ) I48F5E59356CCB45A1C41CAE764DF169C
= I1A7B4E094F07B0C85C5ACADEC807841F ; wire [I20215169A99BAB8B27571CCDC8331264 -1:0] I0F3FCCC5995F6CBAD0568AFF03FA9E41 ; I07DF4961FACFAABF085590F687502283
IC25FB15852E0AA383844DA8C245C8F77 ( .I94A08DA1FECBB6E8B46990538C7B50B2 ({I48F5E59356CCB45A1C41CAE764DF169C , I0F3FCCC5995F6CBAD0568AFF03FA9E41 [I20215169A99BAB8B27571CCDC8331264 -1:1]}),
.ID40B528C645AD71B3CA95E92A7F6C14D (IA70367AA7CB74E510F4F9413CCF059D3 ) ); wire [I20215169A99BAB8B27571CCDC8331264 -1:0]
I8658C20F212661D73D29B60629113469 , IAB790A5ACD86FC696B2B001A6A044D14 , IEA116DC1225420B07D123EB3C08534C0 , I6D43C706A2D0C921C11B984E62071A12 ,
I64D2346B95D903D0423261A186BC883F , IC216F003BDBC623A31E4A8F3AE33C1B1 ; assign I5B9F987DBE3EDAC4E347A14A5782131F
= {I8658C20F212661D73D29B60629113469 [31], I8658C20F212661D73D29B60629113469 [32]}; assign I08C038534302D663980480E37D20BC83
= {IAB790A5ACD86FC696B2B001A6A044D14 [31], IAB790A5ACD86FC696B2B001A6A044D14 [32]}; assign I769454D2A8D191F3E322B7B5DF928B5D
= {IEA116DC1225420B07D123EB3C08534C0 [31], IEA116DC1225420B07D123EB3C08534C0 [32]}; assign I01BDC194686F6DC3F502CFA733822312
= {I6D43C706A2D0C921C11B984E62071A12 [31], I6D43C706A2D0C921C11B984E62071A12 [32]}; assign I87B3D78A5F6FFC46951ED28E772E594D
= {I64D2346B95D903D0423261A186BC883F [31], I64D2346B95D903D0423261A186BC883F [32]}; assign I159859469876028CEA112C7C16B1CAF5
= {IC216F003BDBC623A31E4A8F3AE33C1B1 [31], IC216F003BDBC623A31E4A8F3AE33C1B1 [32]}; wire [I20215169A99BAB8B27571CCDC8331264 *2-1:0]
I5367F16813E8B3314F5C3786E492456F ; assign IAE766072895E2EB8B8716944E133AE63 = I5367F16813E8B3314F5C3786E492456F [I20215169A99BAB8B27571CCDC8331264 *2-1:64]; generate genvar
I8CE4B16B22B58894AA86C421E8759DF3 ; for (I8CE4B16B22B58894AA86C421E8759DF3 =0; I8CE4B16B22B58894AA86C421E8759DF3 <I20215169A99BAB8B27571CCDC8331264 ;
I8CE4B16B22B58894AA86C421E8759DF3 =I8CE4B16B22B58894AA86C421E8759DF3 +1) begin : IBC937D9A13D072E24154E92A7A8AD4EF IB51AA32163492596ADA06B22A9206E8F
I57E3E2F56972AC048D6F35E5F0E3AD1E ( .I0A3BC2148686F2B562665C3891507E35 (I0A3BC2148686F2B562665C3891507E35 ), .I86266EE937D97F812A8E57D22B62EE29 (I86266EE937D97F812A8E57D22B62EE29 ), .I27E9DD9482B253AA850544215471D9D5 (I27E9DD9482B253AA850544215471D9D5 ), .IE9DED2DF97E91174FD62E40E248B137D (IE9DED2DF97E91174FD62E40E248B137D ), .I8715FEDE1A202C700CD025C90F3B2421 (I8715FEDE1A202C700CD025C90F3B2421 ), .I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 (I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 ),
.IFC240E6D824E08568AA642A34947FEBC (ICE7D06150E11255C4F8EE2384429A32A [I8CE4B16B22B58894AA86C421E8759DF3 ]), .I5844CE4E8F912137CD0A723AA7A4EBB2 (ICE7D06150E11255C4F8EE2384429A32A [I8CE4B16B22B58894AA86C421E8759DF3 +1]),
.IF7F7CFDB9A31998C4AEFDC5C8BD5937A (IC9A7CC4AB393A8BD2AE6914033F0530B [I8CE4B16B22B58894AA86C421E8759DF3 *2+1:I8CE4B16B22B58894AA86C421E8759DF3 *2]),
.IC68BD984558E67927B382A860837C32F (ID78F9120B5CAEC4D064AF1B7C0EFA923 [I8CE4B16B22B58894AA86C421E8759DF3 *2+1:I8CE4B16B22B58894AA86C421E8759DF3 *2]),
.I47FE879774A01F989D46EFF34BCF4D44 (IF8DEC8403A8BD60501F344A464CBF9AC [I8CE4B16B22B58894AA86C421E8759DF3 ]), .I1A7B4E094F07B0C85C5ACADEC807841F (IF8DEC8403A8BD60501F344A464CBF9AC [I8CE4B16B22B58894AA86C421E8759DF3 +1]), .I0F3FCCC5995F6CBAD0568AFF03FA9E41 (I0F3FCCC5995F6CBAD0568AFF03FA9E41 [I8CE4B16B22B58894AA86C421E8759DF3 ]),
.I082A499B7DDEF3C7897AB842B431A8AD (I082A499B7DDEF3C7897AB842B431A8AD ), .I89C5B8F33C91378743762C771A89F8C4 (I89C5B8F33C91378743762C771A89F8C4 ), .I8357B924AEFCA0FDD29AADC1ABE078FF (I8357B924AEFCA0FDD29AADC1ABE078FF ),
.I21345BCEA5A3A0213882E3493F7CE8A2 (I21345BCEA5A3A0213882E3493F7CE8A2 ), .IE8F9438C61FEFC48890126E846737803 (IE8F9438C61FEFC48890126E846737803 ),
.I00D170E901FDFA8C4D428ECAC839A4AB (I00D170E901FDFA8C4D428ECAC839A4AB ), .I453DD3088EE862556BDD0F58B390F41F (I453DD3088EE862556BDD0F58B390F41F ),
.I182E80B21C5A5F086FE70D9A01554365 (I182E80B21C5A5F086FE70D9A01554365 ), .I346A81471C889B6C72A88423EB28B21A (I346A81471C889B6C72A88423EB28B21A ),
.I0EB8CC186C9B38B7FB99E477EE981265 (I0EB8CC186C9B38B7FB99E477EE981265 ), .IF41F5F2D34464C2F1512CE4A38EAD286 (IF41F5F2D34464C2F1512CE4A38EAD286 ),
.I75D612F1AEBBE1DC3FC1AC2ED5C21E7F (I75D612F1AEBBE1DC3FC1AC2ED5C21E7F ), .IA882574F5206B0DBAB0B61BA8B369A15 (IE22428CCF96CDA9674A939C209AD1000 [I8CE4B16B22B58894AA86C421E8759DF3 ]),
.IE78AFF6FF490ECAC5AFE4B8DF2BDC999 (IE22428CCF96CDA9674A939C209AD1000 [I8CE4B16B22B58894AA86C421E8759DF3 +1]), .I24D24CDA7F2D8B539E4F5C420BD826D9 (I48A355561F0628CB2813BD54EADAA46C [I8CE4B16B22B58894AA86C421E8759DF3 ]), .I61BAAAAF32AC5A7B6FFEBFC244A2D739 (I61BAAAAF32AC5A7B6FFEBFC244A2D739 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I6E03B4F12533CBA29903F1C9DD1E5C3D (I6E03B4F12533CBA29903F1C9DD1E5C3D [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.IAB9D6A507309488CCF13DB3F67F81B63 (IAB9D6A507309488CCF13DB3F67F81B63 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I83FCEFDFE9F9D1C28AB321626447799F (I83FCEFDFE9F9D1C28AB321626447799F [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I1905DD05FA116073F500B593198EED1C (I1905DD05FA116073F500B593198EED1C [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I61E6EBA71A6BFA5A8FE92AB8FABECBBC (I61E6EBA71A6BFA5A8FE92AB8FABECBBC [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I79EB40C7CC07F0A913BA2E8F9D56D33B (I79EB40C7CC07F0A913BA2E8F9D56D33B [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I973092C325E8C2AE92FFF50B0288E777 (I973092C325E8C2AE92FFF50B0288E777 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.IB9445BEC437AE377554E2723C22C52B2 (IB9445BEC437AE377554E2723C22C52B2 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I6A45CBE320E935B06BB0F08ECF1179D4 (I6A45CBE320E935B06BB0F08ECF1179D4 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I0EE48206D3023D05A5AA46FD33711C98 (I0EE48206D3023D05A5AA46FD33711C98 [I8CE4B16B22B58894AA86C421E8759DF3 /32]), .I81414FA30C7BC73A9A778574097A714B (I81414FA30C7BC73A9A778574097A714B [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I4C39D6D4449338A7DA014742DE16FD46 (I4C39D6D4449338A7DA014742DE16FD46 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.ID8E8746A568679217650DF444D98F91E (ID8E8746A568679217650DF444D98F91E [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I30CD5687FB19DAD9CFD43FE994021B00 (I30CD5687FB19DAD9CFD43FE994021B00 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I018477AF087A1484F83E54C386C2EF07 (I018477AF087A1484F83E54C386C2EF07 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I6970ADE3C1C5CEF4BF2ADF425B8B73CB (I6970ADE3C1C5CEF4BF2ADF425B8B73CB [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I4021D2C4A029457D9671036AF92F0AB8 (I4021D2C4A029457D9671036AF92F0AB8 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I6ABED3933223BDB35402C9F56973AB09 (I6ABED3933223BDB35402C9F56973AB09 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I371CC04BDE216A35CEFED5553951955B (I371CC04BDE216A35CEFED5553951955B [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I032B17AEE0B7BC21B073F5A5AF886D30 (I032B17AEE0B7BC21B073F5A5AF886D30 [I8CE4B16B22B58894AA86C421E8759DF3 /32]),
.I64571D3B8AD6548BEF3F326B0C79154D (I64571D3B8AD6548BEF3F326B0C79154D [I8CE4B16B22B58894AA86C421E8759DF3 /32]), .I528FBBEA2163A7F08F8CE87A6486A505 (I8658C20F212661D73D29B60629113469 [I8CE4B16B22B58894AA86C421E8759DF3 ]),
.IFD2E2FBE657226AA9EB0B69C70CEDAF0 (IAB790A5ACD86FC696B2B001A6A044D14 [I8CE4B16B22B58894AA86C421E8759DF3 ]), .I6034EE230C5F2EA0D0828112861916C6 (IEA116DC1225420B07D123EB3C08534C0 [I8CE4B16B22B58894AA86C421E8759DF3 ]),
.I7E211F728072FEA639172DFD7FC475D2 (I6D43C706A2D0C921C11B984E62071A12 [I8CE4B16B22B58894AA86C421E8759DF3 ]), .I4D5E955D6CD9D5E25ED4CE64CF4DC635 (I64D2346B95D903D0423261A186BC883F [I8CE4B16B22B58894AA86C421E8759DF3 ]),
.I94F01074D91205FEBB9204892C80718F (IC216F003BDBC623A31E4A8F3AE33C1B1 [I8CE4B16B22B58894AA86C421E8759DF3 ]), .IAE766072895E2EB8B8716944E133AE63 (I5367F16813E8B3314F5C3786E492456F [I8CE4B16B22B58894AA86C421E8759DF3 *2+1:I8CE4B16B22B58894AA86C421E8759DF3 *2]) ); end
endgenerate endmodule module I39607C0DCC66F95CC21E6ACF9889D96F (I0A3BC2148686F2B562665C3891507E35 , IF927D8348D0B86E1E1452C2EEF729055 ,
IC68271A63DDBC431C307BEB7D2918275 , IEC4D1EB36B22D19728E9D1D23CA84D1C ); input wire I0A3BC2148686F2B562665C3891507E35 ,
IF927D8348D0B86E1E1452C2EEF729055 ; output reg IC68271A63DDBC431C307BEB7D2918275 ; output wire IEC4D1EB36B22D19728E9D1D23CA84D1C ; wire
[3:0] I2817F701D5E1A1181E657251363295FD ; reg [2:0][3:0] I63372A266D42706F4A794AA5AA935E80 ; initial I63372A266D42706F4A794AA5AA935E80
= 0; always @(posedge I0A3BC2148686F2B562665C3891507E35 ) if (IF927D8348D0B86E1E1452C2EEF729055 ==1 && I2817F701D5E1A1181E657251363295FD
== 9) I63372A266D42706F4A794AA5AA935E80 <= {3{4'b0000}}; else if (IF927D8348D0B86E1E1452C2EEF729055 ==0 && I2817F701D5E1A1181E657251363295FD
== 7) I63372A266D42706F4A794AA5AA935E80 <= {3{4'b0000}}; else I63372A266D42706F4A794AA5AA935E80 <= {3{4'(I2817F701D5E1A1181E657251363295FD +1)}}; assign
I2817F701D5E1A1181E657251363295FD = ( ( I63372A266D42706F4A794AA5AA935E80 [0] & I63372A266D42706F4A794AA5AA935E80 [1]
) | ( I63372A266D42706F4A794AA5AA935E80 [1] & I63372A266D42706F4A794AA5AA935E80 [2] ) | ( I63372A266D42706F4A794AA5AA935E80 [0]
& I63372A266D42706F4A794AA5AA935E80 [2] ) ); always @(posedge I0A3BC2148686F2B562665C3891507E35 ) IC68271A63DDBC431C307BEB7D2918275
<= I2817F701D5E1A1181E657251363295FD [2]; wire I3F76FA0DD412AED50E4391D2F1A23AE3 ; assign I3F76FA0DD412AED50E4391D2F1A23AE3
= (I2817F701D5E1A1181E657251363295FD == 3); reg [2:0] I9FE3A3FED1E89843DF8CCA8C22443856 ; always @(posedge I0A3BC2148686F2B562665C3891507E35 ) I9FE3A3FED1E89843DF8CCA8C22443856
<= {3{I3F76FA0DD412AED50E4391D2F1A23AE3 }}; assign IEC4D1EB36B22D19728E9D1D23CA84D1C = ( ( I9FE3A3FED1E89843DF8CCA8C22443856 [0]
& I9FE3A3FED1E89843DF8CCA8C22443856 [1] ) | ( I9FE3A3FED1E89843DF8CCA8C22443856 [1] & I9FE3A3FED1E89843DF8CCA8C22443856 [2]
) | ( I9FE3A3FED1E89843DF8CCA8C22443856 [0] & I9FE3A3FED1E89843DF8CCA8C22443856 [2] ) ); endmodule module I84F6FB7CD5CD53B5679489A29396448F (I0A3BC2148686F2B562665C3891507E35 ,
IEC4D1EB36B22D19728E9D1D23CA84D1C , I13B5BFE96F3E2FE411C9F66F4A582ADF , IC68271A63DDBC431C307BEB7D2918275 ); input
wire I0A3BC2148686F2B562665C3891507E35 , IEC4D1EB36B22D19728E9D1D23CA84D1C ; input wire [9:0] I13B5BFE96F3E2FE411C9F66F4A582ADF ; output
wire IC68271A63DDBC431C307BEB7D2918275 ; reg [9:0] I2AB64F4EE279E5BAF7AB7059B15E6D12 ; reg [2:0][9:0] IE07BBFCDCAA6E02C3FD7417636615CF7 ; always
@(posedge I0A3BC2148686F2B562665C3891507E35 ) if (IEC4D1EB36B22D19728E9D1D23CA84D1C ) IE07BBFCDCAA6E02C3FD7417636615CF7
<= {3{I13B5BFE96F3E2FE411C9F66F4A582ADF }}; else IE07BBFCDCAA6E02C3FD7417636615CF7 <= {3{I2AB64F4EE279E5BAF7AB7059B15E6D12 [8:0],
1'b0}}; assign I2AB64F4EE279E5BAF7AB7059B15E6D12 = ( ( IE07BBFCDCAA6E02C3FD7417636615CF7 [0] & IE07BBFCDCAA6E02C3FD7417636615CF7 [1]
) | ( IE07BBFCDCAA6E02C3FD7417636615CF7 [1] & IE07BBFCDCAA6E02C3FD7417636615CF7 [2] ) | ( IE07BBFCDCAA6E02C3FD7417636615CF7 [0]
& IE07BBFCDCAA6E02C3FD7417636615CF7 [2] ) ); assign IC68271A63DDBC431C307BEB7D2918275 = I2AB64F4EE279E5BAF7AB7059B15E6D12 [9]; endmodule module
I67D38CAA7C80960859CB2AFCF45A4106 ( input logic I86266EE937D97F812A8E57D22B62EE29 , I0A3BC2148686F2B562665C3891507E35 ,
IF698F67F5666AFF10729D8A1CB1C14D2 , input logic I459A6F79AD9B13CBCB5F692D2CC7A94D , IE7D31FC0602FB2EDE144D18CDFFD816B , output
logic I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 , I2C0F741D5E54A03052A7BAEB8CEFA690 , output logic [3:0] I43938353D4FB12C9720D1A7A7537E069 ,
I6413911CE482DB3AB245D5F066541602 , output wire [23:0] IE55603E44DA0CE59B3E8963A06AA6E5A , output wire ICB7658367C9FDD7110EBE09C34077D2C ,
I2AE05249E15E8C6BF7F6AB2A4306FACA , IC68AD92486D949E2FF7EE4E70CD71E8E ); wire I860D2181FADACEB00A90FAFE2CE53F2C ; assign
I860D2181FADACEB00A90FAFE2CE53F2C = I0A3BC2148686F2B562665C3891507E35 ; localparam I2C070FADF478427A55F05FC54FA9BDA2
= 2; enum {I29D21D89F14D787007DB8BED4B086C3D , ID935F4BB38160520D3CBE34D746068C9 , ICCB2642CF9695C335A736FE838BC2674 ,
IA0206CB0A7A680F7E469BCAE562AF789 , I3466FAB4975481651940ED328AA990E4 } I9ED39E2EA931586B6A985A6942EF573E , I5C65729C8776677E9E07C1FB58B7468C ; always @(posedge
I860D2181FADACEB00A90FAFE2CE53F2C ) if (I86266EE937D97F812A8E57D22B62EE29 ) I9ED39E2EA931586B6A985A6942EF573E <=
I29D21D89F14D787007DB8BED4B086C3D ; else I9ED39E2EA931586B6A985A6942EF573E <= I5C65729C8776677E9E07C1FB58B7468C ; logic
[2:0] I3BD5379BC1D1857D75CBB011DE605466 ; logic [3:0] I7151179D6DF8F1902B355FF2B07829AE , I3666B81AB7FC8B4F62E26BA6FB5C11CB ; logic
I0BDAEE649E8C88C7CE90631AF04B4A34 ; always @(*) begin : ICD5B5F7D68F72B5A6A8AF6EC47E5D5AE I5C65729C8776677E9E07C1FB58B7468C
= I9ED39E2EA931586B6A985A6942EF573E ; case (I9ED39E2EA931586B6A985A6942EF573E ) I29D21D89F14D787007DB8BED4B086C3D
: if (I0BDAEE649E8C88C7CE90631AF04B4A34 ) I5C65729C8776677E9E07C1FB58B7468C = ID935F4BB38160520D3CBE34D746068C9 ;
ID935F4BB38160520D3CBE34D746068C9 : I5C65729C8776677E9E07C1FB58B7468C = ICCB2642CF9695C335A736FE838BC2674 ; ICCB2642CF9695C335A736FE838BC2674
: if (I3BD5379BC1D1857D75CBB011DE605466 == I2C070FADF478427A55F05FC54FA9BDA2 & IE7D31FC0602FB2EDE144D18CDFFD816B
== 1) begin if (I459A6F79AD9B13CBCB5F692D2CC7A94D ) I5C65729C8776677E9E07C1FB58B7468C = IA0206CB0A7A680F7E469BCAE562AF789 ; else
if (I3666B81AB7FC8B4F62E26BA6FB5C11CB != I7151179D6DF8F1902B355FF2B07829AE ) I5C65729C8776677E9E07C1FB58B7468C =
ID935F4BB38160520D3CBE34D746068C9 ; else I5C65729C8776677E9E07C1FB58B7468C = I29D21D89F14D787007DB8BED4B086C3D ; end IA0206CB0A7A680F7E469BCAE562AF789
: I5C65729C8776677E9E07C1FB58B7468C = I3466FAB4975481651940ED328AA990E4 ; I3466FAB4975481651940ED328AA990E4 : if (I3BD5379BC1D1857D75CBB011DE605466
== I2C070FADF478427A55F05FC54FA9BDA2 & IE7D31FC0602FB2EDE144D18CDFFD816B == 1) begin if (I459A6F79AD9B13CBCB5F692D2CC7A94D ) I5C65729C8776677E9E07C1FB58B7468C
= IA0206CB0A7A680F7E469BCAE562AF789 ; else if (I3666B81AB7FC8B4F62E26BA6FB5C11CB != I7151179D6DF8F1902B355FF2B07829AE ) I5C65729C8776677E9E07C1FB58B7468C
= ID935F4BB38160520D3CBE34D746068C9 ; else I5C65729C8776677E9E07C1FB58B7468C = I29D21D89F14D787007DB8BED4B086C3D ; end
endcase end always @(posedge I860D2181FADACEB00A90FAFE2CE53F2C ) if (I86266EE937D97F812A8E57D22B62EE29 || (I9ED39E2EA931586B6A985A6942EF573E
== ID935F4BB38160520D3CBE34D746068C9 || I9ED39E2EA931586B6A985A6942EF573E ==IA0206CB0A7A680F7E469BCAE562AF789 )
) I3BD5379BC1D1857D75CBB011DE605466 <= 0; else if ( I3BD5379BC1D1857D75CBB011DE605466 != I2C070FADF478427A55F05FC54FA9BDA2 ) I3BD5379BC1D1857D75CBB011DE605466
<= I3BD5379BC1D1857D75CBB011DE605466 + 1; always @(posedge I860D2181FADACEB00A90FAFE2CE53F2C ) if (I86266EE937D97F812A8E57D22B62EE29 ) #5ns
I7151179D6DF8F1902B355FF2B07829AE <= 0; else if ( I0BDAEE649E8C88C7CE90631AF04B4A34 && I7151179D6DF8F1902B355FF2B07829AE
+1 != I3666B81AB7FC8B4F62E26BA6FB5C11CB ) #5ns I7151179D6DF8F1902B355FF2B07829AE <= I7151179D6DF8F1902B355FF2B07829AE
+ 1; logic IDD60BEEBCBBD2685650352EA033D9494 ; assign IDD60BEEBCBBD2685650352EA033D9494 = (I3666B81AB7FC8B4F62E26BA6FB5C11CB
!= I7151179D6DF8F1902B355FF2B07829AE && !I459A6F79AD9B13CBCB5F692D2CC7A94D ) && (ICB7658367C9FDD7110EBE09C34077D2C
|| (I9ED39E2EA931586B6A985A6942EF573E ==ICCB2642CF9695C335A736FE838BC2674 && I3BD5379BC1D1857D75CBB011DE605466 ==
I2C070FADF478427A55F05FC54FA9BDA2 & IE7D31FC0602FB2EDE144D18CDFFD816B )); always @(posedge I860D2181FADACEB00A90FAFE2CE53F2C ) if (I86266EE937D97F812A8E57D22B62EE29 ) #5ns
I3666B81AB7FC8B4F62E26BA6FB5C11CB <= 0; else if ( IDD60BEEBCBBD2685650352EA033D9494 ) #5ns I3666B81AB7FC8B4F62E26BA6FB5C11CB
<= I3666B81AB7FC8B4F62E26BA6FB5C11CB + 1; assign I43938353D4FB12C9720D1A7A7537E069 = (I7151179D6DF8F1902B355FF2B07829AE
>> 1) ^ I7151179D6DF8F1902B355FF2B07829AE ; assign I6413911CE482DB3AB245D5F066541602 = (I3666B81AB7FC8B4F62E26BA6FB5C11CB
>> 1) ^ I3666B81AB7FC8B4F62E26BA6FB5C11CB ; always @(posedge I860D2181FADACEB00A90FAFE2CE53F2C ) I0BDAEE649E8C88C7CE90631AF04B4A34
<= IF698F67F5666AFF10729D8A1CB1C14D2 ; assign I2C0F741D5E54A03052A7BAEB8CEFA690 = I0BDAEE649E8C88C7CE90631AF04B4A34 ;
logic ICE87C41B76B3D0572202C382CBDB44CD ; always @(posedge I860D2181FADACEB00A90FAFE2CE53F2C ) if (I9ED39E2EA931586B6A985A6942EF573E
== IA0206CB0A7A680F7E469BCAE562AF789 || (I9ED39E2EA931586B6A985A6942EF573E == I3466FAB4975481651940ED328AA990E4
&& !(I3BD5379BC1D1857D75CBB011DE605466 == I2C070FADF478427A55F05FC54FA9BDA2 & IE7D31FC0602FB2EDE144D18CDFFD816B
== 1))) ICE87C41B76B3D0572202C382CBDB44CD <= 1; else ICE87C41B76B3D0572202C382CBDB44CD <= 0; assign I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4
= ICE87C41B76B3D0572202C382CBDB44CD ; assign ICB7658367C9FDD7110EBE09C34077D2C = (I9ED39E2EA931586B6A985A6942EF573E
== I3466FAB4975481651940ED328AA990E4 && I3BD5379BC1D1857D75CBB011DE605466 == I2C070FADF478427A55F05FC54FA9BDA2 &
IE7D31FC0602FB2EDE144D18CDFFD816B ); assign IC68AD92486D949E2FF7EE4E70CD71E8E = (I5C65729C8776677E9E07C1FB58B7468C
== ID935F4BB38160520D3CBE34D746068C9 ); assign I2AE05249E15E8C6BF7F6AB2A4306FACA = (I9ED39E2EA931586B6A985A6942EF573E
== ICCB2642CF9695C335A736FE838BC2674 && I3BD5379BC1D1857D75CBB011DE605466 == I2C070FADF478427A55F05FC54FA9BDA2 &&
IE7D31FC0602FB2EDE144D18CDFFD816B && (I5C65729C8776677E9E07C1FB58B7468C == ID935F4BB38160520D3CBE34D746068C9 ||
I5C65729C8776677E9E07C1FB58B7468C == IA0206CB0A7A680F7E469BCAE562AF789 )); reg [23:0] I5C5CB5B0EEA849C8D311276622E64891 ; always @(posedge
I860D2181FADACEB00A90FAFE2CE53F2C ) if (I86266EE937D97F812A8E57D22B62EE29 ) I5C5CB5B0EEA849C8D311276622E64891 <=
-1; else I5C5CB5B0EEA849C8D311276622E64891 <= I5C5CB5B0EEA849C8D311276622E64891 + 1; reg [23:0] IA05D076258C4FF44BA0995381537AAAF
[15:0]; always @(posedge I860D2181FADACEB00A90FAFE2CE53F2C ) if (I0BDAEE649E8C88C7CE90631AF04B4A34 ) IA05D076258C4FF44BA0995381537AAAF [I7151179D6DF8F1902B355FF2B07829AE ]
<= I5C5CB5B0EEA849C8D311276622E64891 ; assign IE55603E44DA0CE59B3E8963A06AA6E5A = IA05D076258C4FF44BA0995381537AAAF [I3666B81AB7FC8B4F62E26BA6FB5C11CB ]; endmodule
module I6306CEFA3C21256A792AAE49D35F22A1 ( I0A3BC2148686F2B562665C3891507E35 , I86266EE937D97F812A8E57D22B62EE29 ,
I4A5949BC149B714A0BA0BA74394C72F7 , I9EC4C0AFD450CEAC7ADB81C3BCFC9732 , IE9DC924F238FA6CC29465942875FE8F0 , I7C1BDCF7E82A67D7B3F778AF4288BC57 ,
I6E37B4F7E3FEC3FE4C0B18E41D795449 , IECAE13117D6F0584C25A9DA6C8F8415E , IC851AC6DAE2E29984B567E068D572995 , I2B46E1AA6A4A2089A38865C005769980 , I5D66DC68084DBC91ECB34E334C1BC291 , I51E96C20C528EDDF5025F8B0F8448C53 ); input
wire I4A5949BC149B714A0BA0BA74394C72F7 , I9EC4C0AFD450CEAC7ADB81C3BCFC9732 , I0A3BC2148686F2B562665C3891507E35 ,
I86266EE937D97F812A8E57D22B62EE29 , IECAE13117D6F0584C25A9DA6C8F8415E ; input wire [8:0] I5D66DC68084DBC91ECB34E334C1BC291 ,
I51E96C20C528EDDF5025F8B0F8448C53 ; input wire [3:0] IC851AC6DAE2E29984B567E068D572995 ; input wire [3:0] I2B46E1AA6A4A2089A38865C005769980 ; output
reg I7C1BDCF7E82A67D7B3F778AF4288BC57 ; output wire IE9DC924F238FA6CC29465942875FE8F0 ; output wire I6E37B4F7E3FEC3FE4C0B18E41D795449 ; wire
I79905E60B144D2F6C6719B60453DE2AC ; reg IEA2B2676C28C0DB26D39331A336C6B92 ; reg I9F7D0EE82B6A6CA7DDEAE841F3253059 ; reg
[8:0] I886BB73B3156B0AA24AAC99D2DE0B238 ; assign IE9DC924F238FA6CC29465942875FE8F0 = IEA2B2676C28C0DB26D39331A336C6B92
| I9F7D0EE82B6A6CA7DDEAE841F3253059 | I7C1BDCF7E82A67D7B3F778AF4288BC57 ; wire I5CDEE36EF4FFF80C94D5CF936F57C65B ; assign
I79905E60B144D2F6C6719B60453DE2AC = (I886BB73B3156B0AA24AAC99D2DE0B238 ==I51E96C20C528EDDF5025F8B0F8448C53 ) & IEA2B2676C28C0DB26D39331A336C6B92 ;
wire IC9089F3C9ADAF0186F6FFB1EE8D6501C ; I9E18496CBD21D6A02574C0F31F3D3FB7 IB5AB07CDECF9303FF94DB49578282528 (.I6F13D2E1112161FE6F8EA1EDD3F01310 (I0A3BC2148686F2B562665C3891507E35 ),
.I208F156D4A803025C284BB595A7576B4 (I4A5949BC149B714A0BA0BA74394C72F7 | I79905E60B144D2F6C6719B60453DE2AC ), .I3F3B6F139F935CDE0338584380A06130 (IC9089F3C9ADAF0186F6FFB1EE8D6501C ));
always @(negedge IC9089F3C9ADAF0186F6FFB1EE8D6501C ) if (I4A5949BC149B714A0BA0BA74394C72F7 ) I886BB73B3156B0AA24AAC99D2DE0B238
<= I5D66DC68084DBC91ECB34E334C1BC291 ; else I886BB73B3156B0AA24AAC99D2DE0B238 [3:0] <= IC851AC6DAE2E29984B567E068D572995 ;
always @ (posedge IC9089F3C9ADAF0186F6FFB1EE8D6501C or posedge I86266EE937D97F812A8E57D22B62EE29 ) if (I86266EE937D97F812A8E57D22B62EE29 ) IEA2B2676C28C0DB26D39331A336C6B92
<= 0; else if (I4A5949BC149B714A0BA0BA74394C72F7 ) IEA2B2676C28C0DB26D39331A336C6B92 <= 1; else IEA2B2676C28C0DB26D39331A336C6B92
<= 0; wire I83C6B9FFA7CAFB584E170984750AF63E ; assign I83C6B9FFA7CAFB584E170984750AF63E = IECAE13117D6F0584C25A9DA6C8F8415E
| I86266EE937D97F812A8E57D22B62EE29 ; assign I5CDEE36EF4FFF80C94D5CF936F57C65B = !IEA2B2676C28C0DB26D39331A336C6B92
& I9F7D0EE82B6A6CA7DDEAE841F3253059 & ( I886BB73B3156B0AA24AAC99D2DE0B238 [3:0] == I2B46E1AA6A4A2089A38865C005769980
); always @ (negedge IC9089F3C9ADAF0186F6FFB1EE8D6501C or posedge I83C6B9FFA7CAFB584E170984750AF63E ) if (I83C6B9FFA7CAFB584E170984750AF63E ) I9F7D0EE82B6A6CA7DDEAE841F3253059
<= 0; else if (I79905E60B144D2F6C6719B60453DE2AC & I9EC4C0AFD450CEAC7ADB81C3BCFC9732 ) I9F7D0EE82B6A6CA7DDEAE841F3253059
<= 1; assign I6E37B4F7E3FEC3FE4C0B18E41D795449 = I5CDEE36EF4FFF80C94D5CF936F57C65B ; always @(IECAE13117D6F0584C25A9DA6C8F8415E
or I6E37B4F7E3FEC3FE4C0B18E41D795449 ) if ( IECAE13117D6F0584C25A9DA6C8F8415E == 1'b0 ) I7C1BDCF7E82A67D7B3F778AF4288BC57
= I6E37B4F7E3FEC3FE4C0B18E41D795449 ; endmodule module I4A7799F98F8BFA916086832ADA73E798 #(parameter I6DF7E246C71D6D2493823379E5C1AA50
= 34, parameter IDBF04E8E8F1F83557BAE7BEA2CBD57BD = 2) ( output wire [I6DF7E246C71D6D2493823379E5C1AA50 -1:0] I5316F360783B270FE9AC3887CE27EF1D , output
wire IE01D0BDC7D5682BCB747F7EEFBE73DCB , output wire I561AF95BF4F6EB0D6654C5812AB28B1F , input wire [I6DF7E246C71D6D2493823379E5C1AA50 -1:0]
IA776DD7EA52A4C6B834F3E481B7BDC1F , input wire I72A3034E1DBCB3283E6B3211A628FBD8 , I9AB96B3F1E8B9326C3C792CB4B2BA759 ,
I5814C91DB64F071BEEAA8913CE4B41D9 , input wire I9B05D4C8F2C4E4DEE91A9C511A75634B , I444A7039B02C6D02C8913AA00CF03207 ,
I480B3FA2D679840798F74A04A6C7C705 ); wire [IDBF04E8E8F1F83557BAE7BEA2CBD57BD -1:0] IF5A6A6543A183EE75B3D301249C00DC2 ,
IECCD98B0F221831ACCE46A7EE6F8D293 ; wire [IDBF04E8E8F1F83557BAE7BEA2CBD57BD :0] IEBAE30206FBDF2853755A4FBB0192D6A ,
I853F1D108FE776C69FE2BAADD813A6A1 , I2FABBFEA0AD45B0886AC66759DED2FC3 , I550C2F1F8114167965699309C119BCB1 ; I607CD3EEDA83BC60F7451AB0336B37E6
#(.I719671112AE8A96230446A276595A365 (IDBF04E8E8F1F83557BAE7BEA2CBD57BD )) IB9508866FC10AB15EBF925ABBC5E8CEE (.I2FABBFEA0AD45B0886AC66759DED2FC3 (I2FABBFEA0AD45B0886AC66759DED2FC3 ),
.I853F1D108FE776C69FE2BAADD813A6A1 (I853F1D108FE776C69FE2BAADD813A6A1 ), .I9AB96B3F1E8B9326C3C792CB4B2BA759 (I9AB96B3F1E8B9326C3C792CB4B2BA759 ),
.I5814C91DB64F071BEEAA8913CE4B41D9 (I5814C91DB64F071BEEAA8913CE4B41D9 )); I3078CD6C31A85FD00C2F018F5B0E23B7 #(.I719671112AE8A96230446A276595A365 (IDBF04E8E8F1F83557BAE7BEA2CBD57BD ))
I4F85E62FCBF4125C1CD718670158C943 (.I550C2F1F8114167965699309C119BCB1 (I550C2F1F8114167965699309C119BCB1 ), .IEBAE30206FBDF2853755A4FBB0192D6A (IEBAE30206FBDF2853755A4FBB0192D6A ), .I444A7039B02C6D02C8913AA00CF03207 (I444A7039B02C6D02C8913AA00CF03207 ),
.I480B3FA2D679840798F74A04A6C7C705 (I480B3FA2D679840798F74A04A6C7C705 )); I98F4B119FEDA52829A8231681C7047E0 #(.I0EBD9CC770F78AB57EB145683A007687 (I6DF7E246C71D6D2493823379E5C1AA50 ),
.I719671112AE8A96230446A276595A365 (IDBF04E8E8F1F83557BAE7BEA2CBD57BD )) I3262F1F086CA619B18BB8B7FD2391F4E (.I5316F360783B270FE9AC3887CE27EF1D (I5316F360783B270FE9AC3887CE27EF1D ),
.IA776DD7EA52A4C6B834F3E481B7BDC1F (IA776DD7EA52A4C6B834F3E481B7BDC1F ), .IF5A6A6543A183EE75B3D301249C00DC2 (IF5A6A6543A183EE75B3D301249C00DC2 ),
.IECCD98B0F221831ACCE46A7EE6F8D293 (IECCD98B0F221831ACCE46A7EE6F8D293 ), .IB8EC7C7B4FE8BCE2CD52A52E649A9696 (I72A3034E1DBCB3283E6B3211A628FBD8 ),
.IE01D0BDC7D5682BCB747F7EEFBE73DCB (IE01D0BDC7D5682BCB747F7EEFBE73DCB ), .I9AB96B3F1E8B9326C3C792CB4B2BA759 (I9AB96B3F1E8B9326C3C792CB4B2BA759 )); I6ADE3FFFCABE5BF8F59751F9FACFA746
#(.I719671112AE8A96230446A276595A365 (IDBF04E8E8F1F83557BAE7BEA2CBD57BD )) IF24393249E67E0BCF67D37F88E07D101 (.I561AF95BF4F6EB0D6654C5812AB28B1F (I561AF95BF4F6EB0D6654C5812AB28B1F ), .IECCD98B0F221831ACCE46A7EE6F8D293 (IECCD98B0F221831ACCE46A7EE6F8D293 ), .I853F1D108FE776C69FE2BAADD813A6A1 (I853F1D108FE776C69FE2BAADD813A6A1 ),
.I550C2F1F8114167965699309C119BCB1 (I550C2F1F8114167965699309C119BCB1 ), .I9B05D4C8F2C4E4DEE91A9C511A75634B (I9B05D4C8F2C4E4DEE91A9C511A75634B ),
.I444A7039B02C6D02C8913AA00CF03207 (I444A7039B02C6D02C8913AA00CF03207 ), .I480B3FA2D679840798F74A04A6C7C705 (I480B3FA2D679840798F74A04A6C7C705 )); I112AC8EFCA406EB602C9D1CD565B9925
#(.I719671112AE8A96230446A276595A365 (IDBF04E8E8F1F83557BAE7BEA2CBD57BD )) I1286D327C34DD798157ABD3BA3B1184A (.IE01D0BDC7D5682BCB747F7EEFBE73DCB (IE01D0BDC7D5682BCB747F7EEFBE73DCB ),
.IF5A6A6543A183EE75B3D301249C00DC2 (IF5A6A6543A183EE75B3D301249C00DC2 ), .IEBAE30206FBDF2853755A4FBB0192D6A (IEBAE30206FBDF2853755A4FBB0192D6A ),
.I2FABBFEA0AD45B0886AC66759DED2FC3 (I2FABBFEA0AD45B0886AC66759DED2FC3 ), .I72A3034E1DBCB3283E6B3211A628FBD8 (I72A3034E1DBCB3283E6B3211A628FBD8 ),
.I9AB96B3F1E8B9326C3C792CB4B2BA759 (I9AB96B3F1E8B9326C3C792CB4B2BA759 ), .I5814C91DB64F071BEEAA8913CE4B41D9 (I5814C91DB64F071BEEAA8913CE4B41D9 )); endmodule module
I98F4B119FEDA52829A8231681C7047E0 #(parameter I0EBD9CC770F78AB57EB145683A007687 = 34, parameter I719671112AE8A96230446A276595A365
= 2) ( output wire [I0EBD9CC770F78AB57EB145683A007687 -1:0] I5316F360783B270FE9AC3887CE27EF1D , input wire [I0EBD9CC770F78AB57EB145683A007687 -1:0]
IA776DD7EA52A4C6B834F3E481B7BDC1F , input wire [I719671112AE8A96230446A276595A365 -1:0] IF5A6A6543A183EE75B3D301249C00DC2 ,
IECCD98B0F221831ACCE46A7EE6F8D293 , input wire IB8EC7C7B4FE8BCE2CD52A52E649A9696 , IE01D0BDC7D5682BCB747F7EEFBE73DCB ,
I9AB96B3F1E8B9326C3C792CB4B2BA759 ); localparam IAA1780B4FCCE2D5D9AF13DC25386D111 = 1<<I719671112AE8A96230446A276595A365 ; reg
[I0EBD9CC770F78AB57EB145683A007687 -1:0] I818B3A7C83EE9C6DA4E7195A1E2887EB [0:IAA1780B4FCCE2D5D9AF13DC25386D111 -1]; assign
I5316F360783B270FE9AC3887CE27EF1D = I818B3A7C83EE9C6DA4E7195A1E2887EB [IECCD98B0F221831ACCE46A7EE6F8D293 ]; always
@(posedge I9AB96B3F1E8B9326C3C792CB4B2BA759 ) if (IB8EC7C7B4FE8BCE2CD52A52E649A9696 && !IE01D0BDC7D5682BCB747F7EEFBE73DCB )
I818B3A7C83EE9C6DA4E7195A1E2887EB [IF5A6A6543A183EE75B3D301249C00DC2 ] <= IA776DD7EA52A4C6B834F3E481B7BDC1F ; endmodule module
I6ADE3FFFCABE5BF8F59751F9FACFA746 #(parameter I719671112AE8A96230446A276595A365 = 2) ( output reg I561AF95BF4F6EB0D6654C5812AB28B1F , output
wire [I719671112AE8A96230446A276595A365 -1:0] IECCD98B0F221831ACCE46A7EE6F8D293 , output reg [I719671112AE8A96230446A276595A365
:0] I853F1D108FE776C69FE2BAADD813A6A1 , input wire [I719671112AE8A96230446A276595A365 :0] I550C2F1F8114167965699309C119BCB1 , input
wire I9B05D4C8F2C4E4DEE91A9C511A75634B , I444A7039B02C6D02C8913AA00CF03207 , I480B3FA2D679840798F74A04A6C7C705 ); reg
[I719671112AE8A96230446A276595A365 :0] I89A167FFFCEDF5ACB5885ABD6EF3D145 ; wire [I719671112AE8A96230446A276595A365 :0]
IE424109D3F7B2708274DAC6558278EC4 , I3A9F204D9195CA2A65932949DE9C02D1 ; always @(posedge I444A7039B02C6D02C8913AA00CF03207 ) if
(I480B3FA2D679840798F74A04A6C7C705 ) {I89A167FFFCEDF5ACB5885ABD6EF3D145 , I853F1D108FE776C69FE2BAADD813A6A1 } <=
0; else {I89A167FFFCEDF5ACB5885ABD6EF3D145 , I853F1D108FE776C69FE2BAADD813A6A1 } <= {I3A9F204D9195CA2A65932949DE9C02D1 ,
IE424109D3F7B2708274DAC6558278EC4 }; assign IECCD98B0F221831ACCE46A7EE6F8D293 = I89A167FFFCEDF5ACB5885ABD6EF3D145 [I719671112AE8A96230446A276595A365 -1:0]; assign
I3A9F204D9195CA2A65932949DE9C02D1 = I89A167FFFCEDF5ACB5885ABD6EF3D145 + (I9B05D4C8F2C4E4DEE91A9C511A75634B & ~I561AF95BF4F6EB0D6654C5812AB28B1F ); assign
IE424109D3F7B2708274DAC6558278EC4 = (I3A9F204D9195CA2A65932949DE9C02D1 >>1) ^ I3A9F204D9195CA2A65932949DE9C02D1 ; wire
IDA7B93E3C8E6FC096AAC165560E32370 ; assign IDA7B93E3C8E6FC096AAC165560E32370 = (IE424109D3F7B2708274DAC6558278EC4
== I550C2F1F8114167965699309C119BCB1 ); always @(posedge I444A7039B02C6D02C8913AA00CF03207 ) if (I480B3FA2D679840798F74A04A6C7C705 )
I561AF95BF4F6EB0D6654C5812AB28B1F <= 1'b1; else I561AF95BF4F6EB0D6654C5812AB28B1F <= IDA7B93E3C8E6FC096AAC165560E32370 ; endmodule module
I112AC8EFCA406EB602C9D1CD565B9925 #(parameter I719671112AE8A96230446A276595A365 = 2) ( output reg IE01D0BDC7D5682BCB747F7EEFBE73DCB , output
wire [I719671112AE8A96230446A276595A365 -1:0] IF5A6A6543A183EE75B3D301249C00DC2 , output reg [I719671112AE8A96230446A276595A365
:0] IEBAE30206FBDF2853755A4FBB0192D6A , input wire [I719671112AE8A96230446A276595A365 :0] I2FABBFEA0AD45B0886AC66759DED2FC3 , input
wire I72A3034E1DBCB3283E6B3211A628FBD8 , I9AB96B3F1E8B9326C3C792CB4B2BA759 , I5814C91DB64F071BEEAA8913CE4B41D9 ); reg
[I719671112AE8A96230446A276595A365 :0] IB7DF8095D0F6233307DD8D7D54FE0603 ; wire [I719671112AE8A96230446A276595A365 :0]
IF6714F63E66193A6A6BB65FD5546303A , I89B88BDADF90E6632ABF0632C34E607B ; always @(posedge I9AB96B3F1E8B9326C3C792CB4B2BA759 ) if
(I5814C91DB64F071BEEAA8913CE4B41D9 ) {IB7DF8095D0F6233307DD8D7D54FE0603 , IEBAE30206FBDF2853755A4FBB0192D6A } <=
0; else {IB7DF8095D0F6233307DD8D7D54FE0603 , IEBAE30206FBDF2853755A4FBB0192D6A } <= {I89B88BDADF90E6632ABF0632C34E607B ,
IF6714F63E66193A6A6BB65FD5546303A }; assign IF5A6A6543A183EE75B3D301249C00DC2 = IB7DF8095D0F6233307DD8D7D54FE0603 [I719671112AE8A96230446A276595A365 -1:0]; assign
I89B88BDADF90E6632ABF0632C34E607B = IB7DF8095D0F6233307DD8D7D54FE0603 + (I72A3034E1DBCB3283E6B3211A628FBD8 & ~IE01D0BDC7D5682BCB747F7EEFBE73DCB ); assign
IF6714F63E66193A6A6BB65FD5546303A = (I89B88BDADF90E6632ABF0632C34E607B >>1) ^ I89B88BDADF90E6632ABF0632C34E607B ; wire
I435CCBCF6E534CDB343583716D587417 ; assign I435CCBCF6E534CDB343583716D587417 = (IF6714F63E66193A6A6BB65FD5546303A =={~I2FABBFEA0AD45B0886AC66759DED2FC3 [I719671112AE8A96230446A276595A365 :I719671112AE8A96230446A276595A365 -1],
I2FABBFEA0AD45B0886AC66759DED2FC3 [I719671112AE8A96230446A276595A365 -2:0]}); always @(posedge I9AB96B3F1E8B9326C3C792CB4B2BA759 ) if
(I5814C91DB64F071BEEAA8913CE4B41D9 ) IE01D0BDC7D5682BCB747F7EEFBE73DCB <= 1'b0; else IE01D0BDC7D5682BCB747F7EEFBE73DCB
<= I435CCBCF6E534CDB343583716D587417 ; endmodule module I607CD3EEDA83BC60F7451AB0336B37E6 #(parameter I719671112AE8A96230446A276595A365
= 2) (output reg [I719671112AE8A96230446A276595A365 :0] I2FABBFEA0AD45B0886AC66759DED2FC3 , input wire [I719671112AE8A96230446A276595A365 :0]
I853F1D108FE776C69FE2BAADD813A6A1 , input wire I9AB96B3F1E8B9326C3C792CB4B2BA759 , I5814C91DB64F071BEEAA8913CE4B41D9 ); reg
[I719671112AE8A96230446A276595A365 :0] IF6D130D75AF0CDB6B1BD90FC6C189B20 ; always @(posedge I9AB96B3F1E8B9326C3C792CB4B2BA759 ) if
(I5814C91DB64F071BEEAA8913CE4B41D9 ) {I2FABBFEA0AD45B0886AC66759DED2FC3 ,IF6D130D75AF0CDB6B1BD90FC6C189B20 } <=
0; else {I2FABBFEA0AD45B0886AC66759DED2FC3 ,IF6D130D75AF0CDB6B1BD90FC6C189B20 } <= {IF6D130D75AF0CDB6B1BD90FC6C189B20 ,I853F1D108FE776C69FE2BAADD813A6A1 }; endmodule module
I3078CD6C31A85FD00C2F018F5B0E23B7 #(parameter I719671112AE8A96230446A276595A365 = 2) ( output reg [I719671112AE8A96230446A276595A365 :0]
I550C2F1F8114167965699309C119BCB1 , input wire [I719671112AE8A96230446A276595A365 :0] IEBAE30206FBDF2853755A4FBB0192D6A , input
wire I444A7039B02C6D02C8913AA00CF03207 , I480B3FA2D679840798F74A04A6C7C705 ); reg [I719671112AE8A96230446A276595A365 :0]
I6751318DE9D9D2A14C7FB28D01C6B36F ; always @(posedge I444A7039B02C6D02C8913AA00CF03207 ) if (I480B3FA2D679840798F74A04A6C7C705 )
{I550C2F1F8114167965699309C119BCB1 ,I6751318DE9D9D2A14C7FB28D01C6B36F } <= 0; else {I550C2F1F8114167965699309C119BCB1 ,I6751318DE9D9D2A14C7FB28D01C6B36F }
<= {I6751318DE9D9D2A14C7FB28D01C6B36F ,IEBAE30206FBDF2853755A4FBB0192D6A }; endmodule module I07DF4961FACFAABF085590F687502283 (input
wire [0:63] I94A08DA1FECBB6E8B46990538C7B50B2 , output wire [5:0] ID40B528C645AD71B3CA95E92A7F6C14D ); wire [64:0]
I6EF5B8E14F85B79EA0C56E78FDD4779E [5:0]; generate genvar I8CE4B16B22B58894AA86C421E8759DF3 ; for (I8CE4B16B22B58894AA86C421E8759DF3 =0;
I8CE4B16B22B58894AA86C421E8759DF3 <64; I8CE4B16B22B58894AA86C421E8759DF3 =I8CE4B16B22B58894AA86C421E8759DF3 +1) begin :
I0C9CF0D9833FA8B20E950CB69671BB84 assign I6EF5B8E14F85B79EA0C56E78FDD4779E [0][I8CE4B16B22B58894AA86C421E8759DF3 ]
= !(I6EF5B8E14F85B79EA0C56E78FDD4779E [0][I8CE4B16B22B58894AA86C421E8759DF3 +1] & I94A08DA1FECBB6E8B46990538C7B50B2 [I8CE4B16B22B58894AA86C421E8759DF3 ]); if (I8CE4B16B22B58894AA86C421E8759DF3 %2==0) assign
I6EF5B8E14F85B79EA0C56E78FDD4779E [1][I8CE4B16B22B58894AA86C421E8759DF3 ] = !(I6EF5B8E14F85B79EA0C56E78FDD4779E [1][I8CE4B16B22B58894AA86C421E8759DF3 +2]
& I94A08DA1FECBB6E8B46990538C7B50B2 [I8CE4B16B22B58894AA86C421E8759DF3 ]); if (I8CE4B16B22B58894AA86C421E8759DF3 %4==0) assign
I6EF5B8E14F85B79EA0C56E78FDD4779E [2][I8CE4B16B22B58894AA86C421E8759DF3 ] = !(I6EF5B8E14F85B79EA0C56E78FDD4779E [2][I8CE4B16B22B58894AA86C421E8759DF3 +4]
& I94A08DA1FECBB6E8B46990538C7B50B2 [I8CE4B16B22B58894AA86C421E8759DF3 ]); if (I8CE4B16B22B58894AA86C421E8759DF3 %8==0) assign
I6EF5B8E14F85B79EA0C56E78FDD4779E [3][I8CE4B16B22B58894AA86C421E8759DF3 ] = !(I6EF5B8E14F85B79EA0C56E78FDD4779E [3][I8CE4B16B22B58894AA86C421E8759DF3 +8]
& I94A08DA1FECBB6E8B46990538C7B50B2 [I8CE4B16B22B58894AA86C421E8759DF3 ]); if (I8CE4B16B22B58894AA86C421E8759DF3 %16==0) assign
I6EF5B8E14F85B79EA0C56E78FDD4779E [4][I8CE4B16B22B58894AA86C421E8759DF3 ] = !(I6EF5B8E14F85B79EA0C56E78FDD4779E [4][I8CE4B16B22B58894AA86C421E8759DF3 +16]
& I94A08DA1FECBB6E8B46990538C7B50B2 [I8CE4B16B22B58894AA86C421E8759DF3 ]); if (I8CE4B16B22B58894AA86C421E8759DF3 %32==0) assign
I6EF5B8E14F85B79EA0C56E78FDD4779E [5][I8CE4B16B22B58894AA86C421E8759DF3 ] = !(I6EF5B8E14F85B79EA0C56E78FDD4779E [5][I8CE4B16B22B58894AA86C421E8759DF3 +32]
& I94A08DA1FECBB6E8B46990538C7B50B2 [I8CE4B16B22B58894AA86C421E8759DF3 ]); end endgenerate assign I6EF5B8E14F85B79EA0C56E78FDD4779E [0][64]
= 1; assign I6EF5B8E14F85B79EA0C56E78FDD4779E [1][64] = 1; assign I6EF5B8E14F85B79EA0C56E78FDD4779E [2][64] = 1; assign
I6EF5B8E14F85B79EA0C56E78FDD4779E [3][64] = 1; assign I6EF5B8E14F85B79EA0C56E78FDD4779E [4][64] = 1; assign I6EF5B8E14F85B79EA0C56E78FDD4779E [5][64]
= 1; assign ID40B528C645AD71B3CA95E92A7F6C14D [0] = !I6EF5B8E14F85B79EA0C56E78FDD4779E [0][0]; assign ID40B528C645AD71B3CA95E92A7F6C14D [1]
= !I6EF5B8E14F85B79EA0C56E78FDD4779E [1][0]; assign ID40B528C645AD71B3CA95E92A7F6C14D [2] = !I6EF5B8E14F85B79EA0C56E78FDD4779E [2][0]; assign
ID40B528C645AD71B3CA95E92A7F6C14D [3] = !I6EF5B8E14F85B79EA0C56E78FDD4779E [3][0]; assign ID40B528C645AD71B3CA95E92A7F6C14D [4]
= !I6EF5B8E14F85B79EA0C56E78FDD4779E [4][0]; assign ID40B528C645AD71B3CA95E92A7F6C14D [5] = !I6EF5B8E14F85B79EA0C56E78FDD4779E [5][0]; endmodule
module I89B5FE0A834B8CEFBAD7FEA7A3D23364 ( input IF41F5F2D34464C2F1512CE4A38EAD286 , I75D612F1AEBBE1DC3FC1AC2ED5C21E7F ,
IA882574F5206B0DBAB0B61BA8B369A15 , I0EB8CC186C9B38B7FB99E477EE981265 , output reg IE78AFF6FF490ECAC5AFE4B8DF2BDC999 , input
wire I21345BCEA5A3A0213882E3493F7CE8A2 , input I00D170E901FDFA8C4D428ECAC839A4AB , IE8F9438C61FEFC48890126E846737803 , input
wire [3:0] I182E80B21C5A5F086FE70D9A01554365 , input wire [1:0] I453DD3088EE862556BDD0F58B390F41F , input I346A81471C889B6C72A88423EB28B21A , input
wire IABEB1D6F727D4016CBA8D230E06173E2 , output wire IF365BCF55686BCCD839FE1624DD7D486 , I5FBB67CECBAEE3FB61298BB458246F95 ,
output wire [3:0] IDF6B1552FD717A0BD463ABC2AE6BE59A , I10F9F36D10F50952745A860C2309B5EB , output wire I9415662DEE73FC21C95CE7FCC2E8169E ,
I24D24CDA7F2D8B539E4F5C420BD826D9 ); wire [1:0] I4B2FBF7F994ECB6BD58FA8FB93C5ABF8 ; wire [3:0] I5D3B991ABBF680C2795BD2457E606A8C ; wire
I31C6B3FDFAAA80DBA2DBF92A4600524C ; wire I1E32FC14226F0DBAADFC34BAE0918585 ; reg I943C0B7B2E31ECDE607EC65CC63B9024 ,
I6B9591E70869BF4262EB8D86D58EA914 , I83158F45621E4868B57C91D0579DD86D ; always @(*) begin if (I4B2FBF7F994ECB6BD58FA8FB93C5ABF8
== 2'b00) begin I943C0B7B2E31ECDE607EC65CC63B9024 = 0; I6B9591E70869BF4262EB8D86D58EA914 = 0; I83158F45621E4868B57C91D0579DD86D
= 0; end else if (I4B2FBF7F994ECB6BD58FA8FB93C5ABF8 == 2'b01) begin I943C0B7B2E31ECDE607EC65CC63B9024 = 0; I6B9591E70869BF4262EB8D86D58EA914
= 0; I83158F45621E4868B57C91D0579DD86D = 1; end else if (I4B2FBF7F994ECB6BD58FA8FB93C5ABF8 == 2'b10) begin I943C0B7B2E31ECDE607EC65CC63B9024
= 0; I6B9591E70869BF4262EB8D86D58EA914 = 1; I83158F45621E4868B57C91D0579DD86D = 1; end else begin I943C0B7B2E31ECDE607EC65CC63B9024
= 1; I6B9591E70869BF4262EB8D86D58EA914 = 1; I83158F45621E4868B57C91D0579DD86D = 1; end end reg [1:0] IDD8636B4CE3FEB7420C630CF5F87A588 ; reg
IF40AC107651A7C34D7759E41CBA354C6 , ID74D4F0EC6CE8FE6C2F2A2CA38703336 ; reg [3:0] I2A090335B17F57F393217C6D5EAE3D3F ; always @(*) if (IE8F9438C61FEFC48890126E846737803 ) ID74D4F0EC6CE8FE6C2F2A2CA38703336
= IE78AFF6FF490ECAC5AFE4B8DF2BDC999 ; always @(*) if (I00D170E901FDFA8C4D428ECAC839A4AB ) IF40AC107651A7C34D7759E41CBA354C6
= IE78AFF6FF490ECAC5AFE4B8DF2BDC999 ; generate genvar I8CE4B16B22B58894AA86C421E8759DF3 ; for (I8CE4B16B22B58894AA86C421E8759DF3 =0;
I8CE4B16B22B58894AA86C421E8759DF3 <4; I8CE4B16B22B58894AA86C421E8759DF3 =I8CE4B16B22B58894AA86C421E8759DF3 +1) begin :
I3A94B03CF355E550E11B42CAFDE74D25 always @(*) if (I182E80B21C5A5F086FE70D9A01554365 [I8CE4B16B22B58894AA86C421E8759DF3 ]) I2A090335B17F57F393217C6D5EAE3D3F [I8CE4B16B22B58894AA86C421E8759DF3 ]
= IE78AFF6FF490ECAC5AFE4B8DF2BDC999 ; end endgenerate generate genvar I363B122C528F54DF4A0446B6BAB05515 ; for (I363B122C528F54DF4A0446B6BAB05515 =0;
I363B122C528F54DF4A0446B6BAB05515 <2; I363B122C528F54DF4A0446B6BAB05515 =I363B122C528F54DF4A0446B6BAB05515 +1) begin :
I6885D9C2948C3A01B06CC3ABACF60945 always @(*) if (I453DD3088EE862556BDD0F58B390F41F [I363B122C528F54DF4A0446B6BAB05515 ]) IDD8636B4CE3FEB7420C630CF5F87A588 [I363B122C528F54DF4A0446B6BAB05515 ]
= IE78AFF6FF490ECAC5AFE4B8DF2BDC999 ; end endgenerate wire I550CFD8E2DD2F0382D314AE0EE5CC403 ; assign I550CFD8E2DD2F0382D314AE0EE5CC403
= I75D612F1AEBBE1DC3FC1AC2ED5C21E7F ? IF41F5F2D34464C2F1512CE4A38EAD286 : I9415662DEE73FC21C95CE7FCC2E8169E ; wire
ICEC48D097A13E601ED8E3C25A2BB54DD ; assign ICEC48D097A13E601ED8E3C25A2BB54DD = I75D612F1AEBBE1DC3FC1AC2ED5C21E7F
? IA882574F5206B0DBAB0B61BA8B369A15 : 1'b1; always @(posedge I550CFD8E2DD2F0382D314AE0EE5CC403 ) IE78AFF6FF490ECAC5AFE4B8DF2BDC999
<= ICEC48D097A13E601ED8E3C25A2BB54DD ; assign I4B2FBF7F994ECB6BD58FA8FB93C5ABF8 = I0EB8CC186C9B38B7FB99E477EE981265
? 2'b11 : IDD8636B4CE3FEB7420C630CF5F87A588 ; assign I5FBB67CECBAEE3FB61298BB458246F95 = I0EB8CC186C9B38B7FB99E477EE981265
? 1'b1 : IF40AC107651A7C34D7759E41CBA354C6 ; assign I5D3B991ABBF680C2795BD2457E606A8C = I0EB8CC186C9B38B7FB99E477EE981265
? 4'b1111 : I2A090335B17F57F393217C6D5EAE3D3F ; assign I31C6B3FDFAAA80DBA2DBF92A4600524C = I0EB8CC186C9B38B7FB99E477EE981265
? 1'b0 : ID74D4F0EC6CE8FE6C2F2A2CA38703336 ; assign I1E32FC14226F0DBAADFC34BAE0918585 = I0EB8CC186C9B38B7FB99E477EE981265
? 1'b1 : IE78AFF6FF490ECAC5AFE4B8DF2BDC999 ; wire IEBFE5E1791DB03C4CD6AB95801E0977D ; assign IEBFE5E1791DB03C4CD6AB95801E0977D
= ~IABEB1D6F727D4016CBA8D230E06173E2 ; assign I9415662DEE73FC21C95CE7FCC2E8169E = I21345BCEA5A3A0213882E3493F7CE8A2
? I1E32FC14226F0DBAADFC34BAE0918585 : (IEBFE5E1791DB03C4CD6AB95801E0977D & I6B9591E70869BF4262EB8D86D58EA914 ); assign
I24D24CDA7F2D8B539E4F5C420BD826D9 = I21345BCEA5A3A0213882E3493F7CE8A2 ? I1E32FC14226F0DBAADFC34BAE0918585 : (IEBFE5E1791DB03C4CD6AB95801E0977D
& I943C0B7B2E31ECDE607EC65CC63B9024 ); assign IF365BCF55686BCCD839FE1624DD7D486 = ~I83158F45621E4868B57C91D0579DD86D ; assign
IDF6B1552FD717A0BD463ABC2AE6BE59A = I31C6B3FDFAAA80DBA2DBF92A4600524C ? {4{I346A81471C889B6C72A88423EB28B21A }}
: I5D3B991ABBF680C2795BD2457E606A8C ; assign I10F9F36D10F50952745A860C2309B5EB = I31C6B3FDFAAA80DBA2DBF92A4600524C
? I5D3B991ABBF680C2795BD2457E606A8C : {4{I346A81471C889B6C72A88423EB28B21A }}; endmodule module I9BBBBEA9F740C6E76E42F55F5AB2A5A2
#(parameter I62E5CEF85D46F1A5A2144D9FD463B79E = 1) ( input I0EB8CC186C9B38B7FB99E477EE981265 , I0A3BC2148686F2B562665C3891507E35 ,
I946490AD0FDC17B3B899760A445128F0 , IAC5585D98646D255299C359140537783 , output wire IB807023F87E63B8ADA92F79F546FF9CC , input
[I62E5CEF85D46F1A5A2144D9FD463B79E -1:0] I08804A5B28516A9DC9E56ABFEECF66D9 , output reg [I62E5CEF85D46F1A5A2144D9FD463B79E -1:0]
I7C147CDA9E49590F6ABE83D118B7353B , IE78AFF6FF490ECAC5AFE4B8DF2BDC999 ); always @(posedge I0A3BC2148686F2B562665C3891507E35 ) IE78AFF6FF490ECAC5AFE4B8DF2BDC999
<= {IE78AFF6FF490ECAC5AFE4B8DF2BDC999 [I62E5CEF85D46F1A5A2144D9FD463B79E -2:0], IAC5585D98646D255299C359140537783 }; assign
IB807023F87E63B8ADA92F79F546FF9CC = IE78AFF6FF490ECAC5AFE4B8DF2BDC999 [I62E5CEF85D46F1A5A2144D9FD463B79E -1]; reg
[I62E5CEF85D46F1A5A2144D9FD463B79E -1:0] I8A16ABBC86EBC0B4C2CDAB4364F99F34 ; always @(*) if (I946490AD0FDC17B3B899760A445128F0 ) I8A16ABBC86EBC0B4C2CDAB4364F99F34
= IE78AFF6FF490ECAC5AFE4B8DF2BDC999 ; assign I7C147CDA9E49590F6ABE83D118B7353B = I0EB8CC186C9B38B7FB99E477EE981265
? I08804A5B28516A9DC9E56ABFEECF66D9 : I8A16ABBC86EBC0B4C2CDAB4364F99F34 ; endmodule module IFDB931B30D7BFF08B173BCF1F98E495C (I586A6D64D60A5A9D3DD45E81AA6585A3 ,
I2E192DB878F41E38E0F3B32CFC289D8F , I002953A92DEB31BDFD9E165DFB1DFE1C , I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 , IAE23F82FE849CA57AFF8C2B976AB930E ,
IA5CFBE42922BF86EC0D0DC539D627112 , IFA829BE14FC3FF9B411978DBF7DDF9EE ); parameter I2664F03AC6B8BB9EEE4287720E407DB3
= 1; input wire I586A6D64D60A5A9D3DD45E81AA6585A3 , I2E192DB878F41E38E0F3B32CFC289D8F , I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 ; output
wire I002953A92DEB31BDFD9E165DFB1DFE1C , IAE23F82FE849CA57AFF8C2B976AB930E ; output wire [3:0] IA5CFBE42922BF86EC0D0DC539D627112 ; input
wire [3:0] IFA829BE14FC3FF9B411978DBF7DDF9EE ; assign I002953A92DEB31BDFD9E165DFB1DFE1C = I2E192DB878F41E38E0F3B32CFC289D8F
| I586A6D64D60A5A9D3DD45E81AA6585A3 ; reg I00B57C9FBA005586EC4B8A3796C1E248 ; always @(I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4
or I586A6D64D60A5A9D3DD45E81AA6585A3 ) if (!I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 ) I00B57C9FBA005586EC4B8A3796C1E248
= I586A6D64D60A5A9D3DD45E81AA6585A3 ; reg I68741F9AED41EAAC45E9C8C1AA1F3296 ; always @(I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4
or I2E192DB878F41E38E0F3B32CFC289D8F ) if (!I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 ) I68741F9AED41EAAC45E9C8C1AA1F3296
= I2E192DB878F41E38E0F3B32CFC289D8F ; wire IFE9BCEB45B40932327E66C2EB23FE5ED ; assign IFE9BCEB45B40932327E66C2EB23FE5ED
= (I00B57C9FBA005586EC4B8A3796C1E248 ==0 && I68741F9AED41EAAC45E9C8C1AA1F3296 ==1); wire [3:0] IA18049E0F4D4807E9FD5C8E24DEBD891 ; assign
IA18049E0F4D4807E9FD5C8E24DEBD891 = IFE9BCEB45B40932327E66C2EB23FE5ED ? I2664F03AC6B8BB9EEE4287720E407DB3 : 0; assign
IA5CFBE42922BF86EC0D0DC539D627112 = IA18049E0F4D4807E9FD5C8E24DEBD891 | IFA829BE14FC3FF9B411978DBF7DDF9EE ; assign
IAE23F82FE849CA57AFF8C2B976AB930E = IFE9BCEB45B40932327E66C2EB23FE5ED & I7A1A5F3E79FDC91EDF2F5EAD9D66ABB4 ; endmodule module
I3A7EEC60129C000F5EF89FDB38307204 (ICFE6055D2E0503BE378BB63449EC7BA6 , I9EC4C0AFD450CEAC7ADB81C3BCFC9732 , I86266EE937D97F812A8E57D22B62EE29
,I0A3BC2148686F2B562665C3891507E35 , I47FE879774A01F989D46EFF34BCF4D44 , I1A7B4E094F07B0C85C5ACADEC807841F , IB4CDA117A366592F9BB0BF24B8090648 ,
I662D272D5B777249F5AD3F0BD29F079C , I1653E44E546EA269CD4BEFADAFD0F53C , IC28D2F5880CB3E1E4D819DD6223D52D5 , I37D350E5B2683ED4E78F696D8B080140 ,
IECAE13117D6F0584C25A9DA6C8F8415E , I5EBEE840AC1BD9B012986A05E8BD96CC , I5D66DC68084DBC91ECB34E334C1BC291 , I51E96C20C528EDDF5025F8B0F8448C53 ,
I6F2925832AC361C55FBABB66FC50F914 ); input wire ICFE6055D2E0503BE378BB63449EC7BA6 , I9EC4C0AFD450CEAC7ADB81C3BCFC9732 ,
I86266EE937D97F812A8E57D22B62EE29 , I0A3BC2148686F2B562665C3891507E35 , IB4CDA117A366592F9BB0BF24B8090648 ; input
I6F2925832AC361C55FBABB66FC50F914 ; input wire I47FE879774A01F989D46EFF34BCF4D44 ; output wire I1A7B4E094F07B0C85C5ACADEC807841F ; output
I5EBEE840AC1BD9B012986A05E8BD96CC ; output wire IC28D2F5880CB3E1E4D819DD6223D52D5 ; input wire [3:0] I662D272D5B777249F5AD3F0BD29F079C ; input
wire [3:0] I1653E44E546EA269CD4BEFADAFD0F53C ; output wire [6:0] I37D350E5B2683ED4E78F696D8B080140 ; output wire
[6:0] IECAE13117D6F0584C25A9DA6C8F8415E ; input wire [8:0] I5D66DC68084DBC91ECB34E334C1BC291 , I51E96C20C528EDDF5025F8B0F8448C53 ; wire
[6:0] I7C1BDCF7E82A67D7B3F778AF4288BC57 ; wire [6:0] I6E37B4F7E3FEC3FE4C0B18E41D795449 ; wire [6:0] IE9DC924F238FA6CC29465942875FE8F0 ; wire
[6:0] I07EC8E368A79675BA85B0D28C465226F ; wire [3:0] I8D777F385D3DFEC8815D20F7496026DC [6:0]; generate genvar I8CE4B16B22B58894AA86C421E8759DF3 ; for
(I8CE4B16B22B58894AA86C421E8759DF3 =0; I8CE4B16B22B58894AA86C421E8759DF3 <7; I8CE4B16B22B58894AA86C421E8759DF3 =I8CE4B16B22B58894AA86C421E8759DF3 +1) begin :
IE9A83F5A905606BC889F1E0C5316FC3E I6306CEFA3C21256A792AAE49D35F22A1 IAFC4FC7E48A0710A1DC94EF3E8BC5764 ( .I0A3BC2148686F2B562665C3891507E35 (I0A3BC2148686F2B562665C3891507E35 ),
.I86266EE937D97F812A8E57D22B62EE29 (I86266EE937D97F812A8E57D22B62EE29 ), .I4A5949BC149B714A0BA0BA74394C72F7 (I07EC8E368A79675BA85B0D28C465226F [I8CE4B16B22B58894AA86C421E8759DF3 ]),
.I9EC4C0AFD450CEAC7ADB81C3BCFC9732 (I9EC4C0AFD450CEAC7ADB81C3BCFC9732 ), .IE9DC924F238FA6CC29465942875FE8F0 (IE9DC924F238FA6CC29465942875FE8F0 [I8CE4B16B22B58894AA86C421E8759DF3 ]),
.I7C1BDCF7E82A67D7B3F778AF4288BC57 (I7C1BDCF7E82A67D7B3F778AF4288BC57 [I8CE4B16B22B58894AA86C421E8759DF3 ]), .I6E37B4F7E3FEC3FE4C0B18E41D795449 (I6E37B4F7E3FEC3FE4C0B18E41D795449 [I8CE4B16B22B58894AA86C421E8759DF3 ]),
.IECAE13117D6F0584C25A9DA6C8F8415E (IECAE13117D6F0584C25A9DA6C8F8415E [I8CE4B16B22B58894AA86C421E8759DF3 ]), .IC851AC6DAE2E29984B567E068D572995 (I662D272D5B777249F5AD3F0BD29F079C ),
.I2B46E1AA6A4A2089A38865C005769980 (I1653E44E546EA269CD4BEFADAFD0F53C ), .I5D66DC68084DBC91ECB34E334C1BC291 (I5D66DC68084DBC91ECB34E334C1BC291 ), .I51E96C20C528EDDF5025F8B0F8448C53 (I51E96C20C528EDDF5025F8B0F8448C53 ) ); end
endgenerate wire [6:0] I34E9DC0EA6DE76589A8A1D50E7B0F315 ; generate genvar I6F8F57715090DA2632453988D9A1501B ; for
(I6F8F57715090DA2632453988D9A1501B =0; I6F8F57715090DA2632453988D9A1501B <7; I6F8F57715090DA2632453988D9A1501B =I6F8F57715090DA2632453988D9A1501B +1) begin
: I7B1099C7FF1DDAB1E809FABFF7A7549F if ( I6F8F57715090DA2632453988D9A1501B ==0 ) assign I34E9DC0EA6DE76589A8A1D50E7B0F315 [I6F8F57715090DA2632453988D9A1501B ]
= (IE9DC924F238FA6CC29465942875FE8F0 [I6F8F57715090DA2632453988D9A1501B ]==0); else assign I34E9DC0EA6DE76589A8A1D50E7B0F315 [I6F8F57715090DA2632453988D9A1501B ]
= (IE9DC924F238FA6CC29465942875FE8F0 [I6F8F57715090DA2632453988D9A1501B ]==0 & ( &IE9DC924F238FA6CC29465942875FE8F0 [I6F8F57715090DA2632453988D9A1501B -1:0]
)); end endgenerate assign I07EC8E368A79675BA85B0D28C465226F = {7{ICFE6055D2E0503BE378BB63449EC7BA6 }} & I34E9DC0EA6DE76589A8A1D50E7B0F315
; assign I37D350E5B2683ED4E78F696D8B080140 = I34E9DC0EA6DE76589A8A1D50E7B0F315 ; wire I1A19E3FB6355DFA8D7ACD314EBC49909 ; assign
I1A19E3FB6355DFA8D7ACD314EBC49909 = (I6E37B4F7E3FEC3FE4C0B18E41D795449 != 0); wire I371A650846739DB0C9E8E7A3BA2F181A ;
assign I371A650846739DB0C9E8E7A3BA2F181A = (I1A19E3FB6355DFA8D7ACD314EBC49909 & ~I6F2925832AC361C55FBABB66FC50F914 );
assign I1A7B4E094F07B0C85C5ACADEC807841F = I371A650846739DB0C9E8E7A3BA2F181A | I47FE879774A01F989D46EFF34BCF4D44 ; reg
I48F5E59356CCB45A1C41CAE764DF169C ; always @(I47FE879774A01F989D46EFF34BCF4D44 or IB4CDA117A366592F9BB0BF24B8090648 ) if (
IB4CDA117A366592F9BB0BF24B8090648 == 1'b0 ) I48F5E59356CCB45A1C41CAE764DF169C = I47FE879774A01F989D46EFF34BCF4D44 ; wire
I94035641506BA0549F8B91F84037DE6A ; assign I94035641506BA0549F8B91F84037DE6A = (I48F5E59356CCB45A1C41CAE764DF169C ==0
&& |I7C1BDCF7E82A67D7B3F778AF4288BC57 & IB4CDA117A366592F9BB0BF24B8090648 ); wire [6:0] IEDB71F9ADC72DAEF0301FA4A1B38478E ; generate genvar
IE358EFA489F58062F10DD7316B65649E ; for (IE358EFA489F58062F10DD7316B65649E =0; IE358EFA489F58062F10DD7316B65649E <7;
IE358EFA489F58062F10DD7316B65649E =IE358EFA489F58062F10DD7316B65649E +1) begin : I25501EEA594185D70CDEB6BD9AE5F03C
if ( IE358EFA489F58062F10DD7316B65649E ==0 ) assign IEDB71F9ADC72DAEF0301FA4A1B38478E [IE358EFA489F58062F10DD7316B65649E ]
= (I7C1BDCF7E82A67D7B3F778AF4288BC57 [IE358EFA489F58062F10DD7316B65649E ]==1); else assign IEDB71F9ADC72DAEF0301FA4A1B38478E [IE358EFA489F58062F10DD7316B65649E ]
= (I7C1BDCF7E82A67D7B3F778AF4288BC57 [IE358EFA489F58062F10DD7316B65649E ]==1 & !( |I7C1BDCF7E82A67D7B3F778AF4288BC57 [IE358EFA489F58062F10DD7316B65649E -1:0]
)); end endgenerate assign IECAE13117D6F0584C25A9DA6C8F8415E = I94035641506BA0549F8B91F84037DE6A ? IEDB71F9ADC72DAEF0301FA4A1B38478E
: 0 ; assign IC28D2F5880CB3E1E4D819DD6223D52D5 = I94035641506BA0549F8B91F84037DE6A ; assign I5EBEE840AC1BD9B012986A05E8BD96CC
= I48F5E59356CCB45A1C41CAE764DF169C ; endmodule module IABC6B35F4B0413305137538EE4407E67 (I02F62FEAFD6D93D552D5B8716C48A42B ,
I8CE4B16B22B58894AA86C421E8759DF3 , I1816A803A42A3A548A47FD7B90407CAC , I8F9C634FB2FBC4B39107A845EF6445C6 , I8CD2DE889F491A5FFB5BB3AF153546D5 )
; input [7:0] I02F62FEAFD6D93D552D5B8716C48A42B ; input I8CE4B16B22B58894AA86C421E8759DF3 ; input I1816A803A42A3A548A47FD7B90407CAC
; output [9:0] I8F9C634FB2FBC4B39107A845EF6445C6 ; output I8CD2DE889F491A5FFB5BB3AF153546D5 ; wire I4921C0E2D1F6005ABE1F9EC2E2041909
= I02F62FEAFD6D93D552D5B8716C48A42B [0] ; wire I99D4FB3DB1563C87DA2CDFC0158B37C3 = I02F62FEAFD6D93D552D5B8716C48A42B [1]
; wire I35EA51BAF1FE7F0142AD5F950855DDE0 = I02F62FEAFD6D93D552D5B8716C48A42B [2] ; wire I690382DDCCB8ABC7367A136262E1978F
= I02F62FEAFD6D93D552D5B8716C48A42B [3] ; wire I1EE2225A0118C6A8FF464CF2926CF352 = I02F62FEAFD6D93D552D5B8716C48A42B [4]
; wire I75778BF8FDE7266D416B0089E7B8B793 = I02F62FEAFD6D93D552D5B8716C48A42B [5] ; wire I28DD376C5A44ACC92E450EE338260C56
= I02F62FEAFD6D93D552D5B8716C48A42B [6] ; wire I49F68A5C8493EC2C0BF489821C21FC3B = I02F62FEAFD6D93D552D5B8716C48A42B [7]
; wire I988287F7A1EB966FFC4E19BDBDEEC7C3 = I8CE4B16B22B58894AA86C421E8759DF3 ; wire I85BF921A466C2F6EDA46CFCBE2444D39
= (I4921C0E2D1F6005ABE1F9EC2E2041909 & I99D4FB3DB1563C87DA2CDFC0158B37C3 ) | (!I4921C0E2D1F6005ABE1F9EC2E2041909
& !I99D4FB3DB1563C87DA2CDFC0158B37C3 ) ; wire IEED64930282714BB783BB8650B3F6ED8 = (I35EA51BAF1FE7F0142AD5F950855DDE0
& I690382DDCCB8ABC7367A136262E1978F ) | (!I35EA51BAF1FE7F0142AD5F950855DDE0 & !I690382DDCCB8ABC7367A136262E1978F )
; wire I6A0823D7BC9D11A640A14234F630DA70 = (I4921C0E2D1F6005ABE1F9EC2E2041909 & I99D4FB3DB1563C87DA2CDFC0158B37C3
& !I35EA51BAF1FE7F0142AD5F950855DDE0 & !I690382DDCCB8ABC7367A136262E1978F ) | (I35EA51BAF1FE7F0142AD5F950855DDE0
& I690382DDCCB8ABC7367A136262E1978F & !I4921C0E2D1F6005ABE1F9EC2E2041909 & !I99D4FB3DB1563C87DA2CDFC0158B37C3 )
| ( !I85BF921A466C2F6EDA46CFCBE2444D39 & !IEED64930282714BB783BB8650B3F6ED8 ) ; wire I5CD76C8AF7E804E1F78F03ED85EA3A99
= I4921C0E2D1F6005ABE1F9EC2E2041909 & I99D4FB3DB1563C87DA2CDFC0158B37C3 & I35EA51BAF1FE7F0142AD5F950855DDE0 & I690382DDCCB8ABC7367A136262E1978F
; wire ICC1ED10A86F3A2F553E335032BAD49E3 = !I4921C0E2D1F6005ABE1F9EC2E2041909 & !I99D4FB3DB1563C87DA2CDFC0158B37C3
& !I35EA51BAF1FE7F0142AD5F950855DDE0 & !I690382DDCCB8ABC7367A136262E1978F ; wire I63A9EC78D81D7EB45535FEF90E4012F4
= ( !I85BF921A466C2F6EDA46CFCBE2444D39 & !I35EA51BAF1FE7F0142AD5F950855DDE0 & !I690382DDCCB8ABC7367A136262E1978F )
| ( !IEED64930282714BB783BB8650B3F6ED8 & !I4921C0E2D1F6005ABE1F9EC2E2041909 & !I99D4FB3DB1563C87DA2CDFC0158B37C3 )
; wire I4E6D39E3546BC9B879A80BA506E07B8D = ( !I85BF921A466C2F6EDA46CFCBE2444D39 & I35EA51BAF1FE7F0142AD5F950855DDE0
& I690382DDCCB8ABC7367A136262E1978F ) | ( !IEED64930282714BB783BB8650B3F6ED8 & I4921C0E2D1F6005ABE1F9EC2E2041909
& I99D4FB3DB1563C87DA2CDFC0158B37C3 ) ; wire IADAC5E63F80F8629E9573527B25891D3 = I4921C0E2D1F6005ABE1F9EC2E2041909
; wire IAD7532D5B3860A408FBE01F9455DCA36 = (I99D4FB3DB1563C87DA2CDFC0158B37C3 & !I5CD76C8AF7E804E1F78F03ED85EA3A99 )
| ICC1ED10A86F3A2F553E335032BAD49E3 ; wire IAB6C040066603EF2519D512B21DCE9AB = ICC1ED10A86F3A2F553E335032BAD49E3
| I35EA51BAF1FE7F0142AD5F950855DDE0 | (I1EE2225A0118C6A8FF464CF2926CF352 & I690382DDCCB8ABC7367A136262E1978F & !I35EA51BAF1FE7F0142AD5F950855DDE0
& !I99D4FB3DB1563C87DA2CDFC0158B37C3 & !I4921C0E2D1F6005ABE1F9EC2E2041909 ) ; wire IBF7C782E5C5789716136BC717F227EC5
= I690382DDCCB8ABC7367A136262E1978F & ! (I4921C0E2D1F6005ABE1F9EC2E2041909 & I99D4FB3DB1563C87DA2CDFC0158B37C3 &
I35EA51BAF1FE7F0142AD5F950855DDE0 ) ; wire I504332760740D229CD79CADD87588941 = (I1EE2225A0118C6A8FF464CF2926CF352
| I63A9EC78D81D7EB45535FEF90E4012F4 ) & ! (I1EE2225A0118C6A8FF464CF2926CF352 & I690382DDCCB8ABC7367A136262E1978F
& !I35EA51BAF1FE7F0142AD5F950855DDE0 & !I99D4FB3DB1563C87DA2CDFC0158B37C3 & !I4921C0E2D1F6005ABE1F9EC2E2041909 )
; wire IF98ED07A4D5F50F7DE1410D905F1477F = (I6A0823D7BC9D11A640A14234F630DA70 & !I1EE2225A0118C6A8FF464CF2926CF352 )
| (I1EE2225A0118C6A8FF464CF2926CF352 & !I690382DDCCB8ABC7367A136262E1978F & !I35EA51BAF1FE7F0142AD5F950855DDE0 &
!(I4921C0E2D1F6005ABE1F9EC2E2041909 &I99D4FB3DB1563C87DA2CDFC0158B37C3 )) | (I1EE2225A0118C6A8FF464CF2926CF352 &
I5CD76C8AF7E804E1F78F03ED85EA3A99 ) | (I988287F7A1EB966FFC4E19BDBDEEC7C3 & I1EE2225A0118C6A8FF464CF2926CF352 & I690382DDCCB8ABC7367A136262E1978F
& I35EA51BAF1FE7F0142AD5F950855DDE0 & !I99D4FB3DB1563C87DA2CDFC0158B37C3 & !I4921C0E2D1F6005ABE1F9EC2E2041909 )
| (I1EE2225A0118C6A8FF464CF2926CF352 & !I690382DDCCB8ABC7367A136262E1978F & I35EA51BAF1FE7F0142AD5F950855DDE0 &
!I99D4FB3DB1563C87DA2CDFC0158B37C3 & !I4921C0E2D1F6005ABE1F9EC2E2041909 ) ; wire I714C197AF70D72C2E1911D4E1939C9A9
= (I1EE2225A0118C6A8FF464CF2926CF352 & I690382DDCCB8ABC7367A136262E1978F & !I35EA51BAF1FE7F0142AD5F950855DDE0 &
!I99D4FB3DB1563C87DA2CDFC0158B37C3 & !I4921C0E2D1F6005ABE1F9EC2E2041909 ) | (!I1EE2225A0118C6A8FF464CF2926CF352
& !I6A0823D7BC9D11A640A14234F630DA70 & !I4E6D39E3546BC9B879A80BA506E07B8D ) ; wire I2C605FBD86A134FF29C9BA1ED550BA09
= I988287F7A1EB966FFC4E19BDBDEEC7C3 | (I1EE2225A0118C6A8FF464CF2926CF352 & !I6A0823D7BC9D11A640A14234F630DA70 &
!I63A9EC78D81D7EB45535FEF90E4012F4 ) | (!I1EE2225A0118C6A8FF464CF2926CF352 & !I690382DDCCB8ABC7367A136262E1978F
& I35EA51BAF1FE7F0142AD5F950855DDE0 & I99D4FB3DB1563C87DA2CDFC0158B37C3 & I4921C0E2D1F6005ABE1F9EC2E2041909 ) ; wire
I46C2D303D393C23DF2411CBE2E26574C = I714C197AF70D72C2E1911D4E1939C9A9 ; wire I753B33AD7DB028946F801F3FAF7FC892 =
I988287F7A1EB966FFC4E19BDBDEEC7C3 | (I1EE2225A0118C6A8FF464CF2926CF352 & !I6A0823D7BC9D11A640A14234F630DA70 & !I63A9EC78D81D7EB45535FEF90E4012F4 )
; wire I60C784DE67A671BF846F913183696C05 = I75778BF8FDE7266D416B0089E7B8B793 & I28DD376C5A44ACC92E450EE338260C56
& I49F68A5C8493EC2C0BF489821C21FC3B & (I988287F7A1EB966FFC4E19BDBDEEC7C3 | (I1816A803A42A3A548A47FD7B90407CAC ?
(!I1EE2225A0118C6A8FF464CF2926CF352 & I690382DDCCB8ABC7367A136262E1978F & I4E6D39E3546BC9B879A80BA506E07B8D ) :
(I1EE2225A0118C6A8FF464CF2926CF352 & !I690382DDCCB8ABC7367A136262E1978F & I63A9EC78D81D7EB45535FEF90E4012F4 )))
; wire IEED807024939B808083F0031A56E9872 = I75778BF8FDE7266D416B0089E7B8B793 & ! I60C784DE67A671BF846F913183696C05
; wire I34D1F91FB2E514B8576FAB1A75A89A6B = I28DD376C5A44ACC92E450EE338260C56 | (!I75778BF8FDE7266D416B0089E7B8B793
& !I28DD376C5A44ACC92E450EE338260C56 & !I49F68A5C8493EC2C0BF489821C21FC3B ) ; wire IB5D9B59113086D3F9F9F108ADAAA9AB5
= I49F68A5C8493EC2C0BF489821C21FC3B ; wire I674F33841E2309FFDD24C85DC3B999DE = (!I49F68A5C8493EC2C0BF489821C21FC3B
& (I28DD376C5A44ACC92E450EE338260C56 ^ I75778BF8FDE7266D416B0089E7B8B793 )) | I60C784DE67A671BF846F913183696C05
; wire ID362BAFF82E07002A1FFEC4476672040 = I75778BF8FDE7266D416B0089E7B8B793 & I28DD376C5A44ACC92E450EE338260C56
; wire IAE889B85BB9275E15D7539E53F47CA82 = (!I75778BF8FDE7266D416B0089E7B8B793 & !I28DD376C5A44ACC92E450EE338260C56 )
| (I988287F7A1EB966FFC4E19BDBDEEC7C3 & ((I75778BF8FDE7266D416B0089E7B8B793 & !I28DD376C5A44ACC92E450EE338260C56 )
| (!I75778BF8FDE7266D416B0089E7B8B793 & I28DD376C5A44ACC92E450EE338260C56 ))) ; wire I88881A34CC252F9045E4D8752691489A
= (!I75778BF8FDE7266D416B0089E7B8B793 & !I28DD376C5A44ACC92E450EE338260C56 ) ; wire IBBD6394346DC3136D2FA238A9D3A243D
= I75778BF8FDE7266D416B0089E7B8B793 & I28DD376C5A44ACC92E450EE338260C56 & I49F68A5C8493EC2C0BF489821C21FC3B ; wire
IA71C5C0288C0F345F3666D5F6CA7CA24 = I988287F7A1EB966FFC4E19BDBDEEC7C3 & (I4921C0E2D1F6005ABE1F9EC2E2041909 | I99D4FB3DB1563C87DA2CDFC0158B37C3
| !I35EA51BAF1FE7F0142AD5F950855DDE0 | !I690382DDCCB8ABC7367A136262E1978F | !I1EE2225A0118C6A8FF464CF2926CF352 )
& (!I75778BF8FDE7266D416B0089E7B8B793 | !I28DD376C5A44ACC92E450EE338260C56 | !I49F68A5C8493EC2C0BF489821C21FC3B
| !I1EE2225A0118C6A8FF464CF2926CF352 | !I4E6D39E3546BC9B879A80BA506E07B8D ) ; wire I789CB7C3DCF5D079696EEC4A72C61D76
= (I714C197AF70D72C2E1911D4E1939C9A9 & !I1816A803A42A3A548A47FD7B90407CAC ) | (I2C605FBD86A134FF29C9BA1ED550BA09
& I1816A803A42A3A548A47FD7B90407CAC ) ; wire IF77DDD4D01455C539FB1B57F95B09993 = I1816A803A42A3A548A47FD7B90407CAC
^ (I46C2D303D393C23DF2411CBE2E26574C | I753B33AD7DB028946F801F3FAF7FC892 ) ; wire ID93643F844C740997B9C759ECBB78091
= (IAE889B85BB9275E15D7539E53F47CA82 & !IF77DDD4D01455C539FB1B57F95B09993 ) | (ID362BAFF82E07002A1FFEC4476672040
& IF77DDD4D01455C539FB1B57F95B09993 ) ; assign I8CD2DE889F491A5FFB5BB3AF153546D5 = IF77DDD4D01455C539FB1B57F95B09993
^ (I88881A34CC252F9045E4D8752691489A | IBBD6394346DC3136D2FA238A9D3A243D ) ; assign I8F9C634FB2FBC4B39107A845EF6445C6
= {(I674F33841E2309FFDD24C85DC3B999DE ^ ID93643F844C740997B9C759ECBB78091 ), (IB5D9B59113086D3F9F9F108ADAAA9AB5
^ ID93643F844C740997B9C759ECBB78091 ), (I34D1F91FB2E514B8576FAB1A75A89A6B ^ ID93643F844C740997B9C759ECBB78091 ),
(IEED807024939B808083F0031A56E9872 ^ ID93643F844C740997B9C759ECBB78091 ), (IF98ED07A4D5F50F7DE1410D905F1477F ^ I789CB7C3DCF5D079696EEC4A72C61D76 ),
(I504332760740D229CD79CADD87588941 ^ I789CB7C3DCF5D079696EEC4A72C61D76 ), (IBF7C782E5C5789716136BC717F227EC5 ^ I789CB7C3DCF5D079696EEC4A72C61D76 ),
(IAB6C040066603EF2519D512B21DCE9AB ^ I789CB7C3DCF5D079696EEC4A72C61D76 ), (IAD7532D5B3860A408FBE01F9455DCA36 ^ I789CB7C3DCF5D079696EEC4A72C61D76 ),
(IADAC5E63F80F8629E9573527B25891D3 ^ I789CB7C3DCF5D079696EEC4A72C61D76 )} ; endmodule module I507DE87DD0643D9F2D064D87FF8CE8DD (
input I86266EE937D97F812A8E57D22B62EE29 , I0A3BC2148686F2B562665C3891507E35 , ID9C51D9F54B5E373B300DA2EDDDBB764 , input
[23:0] I8D777F385D3DFEC8815D20F7496026DC , output logic I231E0CDCBF2977BEA26AECDA5A7F45FC , output logic I3D2E8D60C335C528A7C12445BD1F41E3 , output
logic IC68271A63DDBC431C307BEB7D2918275 , input I50BB776CBF75FDBDD857EF107CDA97D3 , input IB4702C9059470087164094C2E5F94070 , input
[7:0] IA55086E1186D1C3CC0FFF510278DF91E , input IB61F32A2FFDFF16751219654FC5AE6E7 ); localparam I1A004F5ABE2B334DB21328BE1EA6B593 =2'b00,
I7AD4905B4543AB4A1637DD23C50E36CE =2'b01 , IE44F9E348E41CB272EFA87387728571B =2'b10, I5C62905D226C50178205CCCDB8C82788 =2'b11; logic
[1:0] I9ED39E2EA931586B6A985A6942EF573E , I5C65729C8776677E9E07C1FB58B7468C ; logic ID5972F1602659028768AC47B9316B673 ; logic
IAD05C732EFA7E73CEB25AFAF7B6B2684 ; assign IAD05C732EFA7E73CEB25AFAF7B6B2684 = !I50BB776CBF75FDBDD857EF107CDA97D3 ; assign
I3D2E8D60C335C528A7C12445BD1F41E3 = ID5972F1602659028768AC47B9316B673 ; logic [1:0] I3EC5B1B4C96DB2313F610F9A4300E221 ; logic
[2:0][1:0] I5941B82B37CEB7CB8E8E8FC9AFAD9701 ; always @(posedge ID5972F1602659028768AC47B9316B673 ) begin if (I86266EE937D97F812A8E57D22B62EE29 ) I5941B82B37CEB7CB8E8E8FC9AFAD9701
<= {3{I1A004F5ABE2B334DB21328BE1EA6B593 }}; else I5941B82B37CEB7CB8E8E8FC9AFAD9701 <= {3{I5C65729C8776677E9E07C1FB58B7468C }}; end assign
I9ED39E2EA931586B6A985A6942EF573E = ( I5941B82B37CEB7CB8E8E8FC9AFAD9701 [0] & I5941B82B37CEB7CB8E8E8FC9AFAD9701 [1]
) | ( I5941B82B37CEB7CB8E8E8FC9AFAD9701 [1] & I5941B82B37CEB7CB8E8E8FC9AFAD9701 [2] ) | ( I5941B82B37CEB7CB8E8E8FC9AFAD9701 [0]
& I5941B82B37CEB7CB8E8E8FC9AFAD9701 [2] ) ; always @(*) begin : ICD5B5F7D68F72B5A6A8AF6EC47E5D5AE I5C65729C8776677E9E07C1FB58B7468C
= I9ED39E2EA931586B6A985A6942EF573E ; case (I9ED39E2EA931586B6A985A6942EF573E ) I1A004F5ABE2B334DB21328BE1EA6B593 : if (ID9C51D9F54B5E373B300DA2EDDDBB764
== 0) I5C65729C8776677E9E07C1FB58B7468C = I7AD4905B4543AB4A1637DD23C50E36CE ; I7AD4905B4543AB4A1637DD23C50E36CE : I5C65729C8776677E9E07C1FB58B7468C
= IE44F9E348E41CB272EFA87387728571B ; IE44F9E348E41CB272EFA87387728571B : if (I3EC5B1B4C96DB2313F610F9A4300E221
== 2) I5C65729C8776677E9E07C1FB58B7468C = I5C62905D226C50178205CCCDB8C82788 ; I5C62905D226C50178205CCCDB8C82788 : if (ID9C51D9F54B5E373B300DA2EDDDBB764
== 1) I5C65729C8776677E9E07C1FB58B7468C = I1A004F5ABE2B334DB21328BE1EA6B593 ; else if (IB61F32A2FFDFF16751219654FC5AE6E7 )
begin if (IAD05C732EFA7E73CEB25AFAF7B6B2684 ) I5C65729C8776677E9E07C1FB58B7468C = I7AD4905B4543AB4A1637DD23C50E36CE ; else
I5C65729C8776677E9E07C1FB58B7468C = I1A004F5ABE2B334DB21328BE1EA6B593 ; end else I5C65729C8776677E9E07C1FB58B7468C
= IE44F9E348E41CB272EFA87387728571B ; endcase end assign I231E0CDCBF2977BEA26AECDA5A7F45FC = ((I9ED39E2EA931586B6A985A6942EF573E
== IE44F9E348E41CB272EFA87387728571B && I3EC5B1B4C96DB2313F610F9A4300E221 == 2)); logic [2:0][1:0] I4179060EE6D7B4132E8F7AE5CAE26254 ; always @(posedge
ID5972F1602659028768AC47B9316B673 ) if (I9ED39E2EA931586B6A985A6942EF573E == I7AD4905B4543AB4A1637DD23C50E36CE ||
I3EC5B1B4C96DB2313F610F9A4300E221 == 2 || I86266EE937D97F812A8E57D22B62EE29 ) I4179060EE6D7B4132E8F7AE5CAE26254
<= {3{2'b00}}; else I4179060EE6D7B4132E8F7AE5CAE26254 <= {3{2'(I3EC5B1B4C96DB2313F610F9A4300E221 + 1)}}; assign
I3EC5B1B4C96DB2313F610F9A4300E221 = ( ( I4179060EE6D7B4132E8F7AE5CAE26254 [0] & I4179060EE6D7B4132E8F7AE5CAE26254 [1]
) | ( I4179060EE6D7B4132E8F7AE5CAE26254 [1] & I4179060EE6D7B4132E8F7AE5CAE26254 [2] ) | ( I4179060EE6D7B4132E8F7AE5CAE26254 [0]
& I4179060EE6D7B4132E8F7AE5CAE26254 [2] ) ); logic [7:0] IE9E97C511899C07C74E75269A2ABA956 ; logic I10315042C15E5BE9C16B02711AC72209 ; logic
I021CFCAE834FA766B3091B6B708D8140 ; logic I363515199821A877761C5143490995BD ; logic [7:0] IB9C5339A9F988BDA02C82F2B8C804151 ; logic
[7:0] IC253D6434FF9417456C113B2B59750EE [2:0]; assign IC253D6434FF9417456C113B2B59750EE [2] = I8D777F385D3DFEC8815D20F7496026DC [7:0];
assign IC253D6434FF9417456C113B2B59750EE [1] = I8D777F385D3DFEC8815D20F7496026DC [15:8]; assign IC253D6434FF9417456C113B2B59750EE [0]
= I8D777F385D3DFEC8815D20F7496026DC [23:16]; logic I93707F725009F066ECF17DD8F6409A66 ; assign I93707F725009F066ECF17DD8F6409A66
= (ID9C51D9F54B5E373B300DA2EDDDBB764 | IB61F32A2FFDFF16751219654FC5AE6E7 ); always @(*) begin if (I9ED39E2EA931586B6A985A6942EF573E
== I7AD4905B4543AB4A1637DD23C50E36CE ) IE9E97C511899C07C74E75269A2ABA956 = 8'b111_11100; else if (I9ED39E2EA931586B6A985A6942EF573E
== IE44F9E348E41CB272EFA87387728571B ) IE9E97C511899C07C74E75269A2ABA956 = IC253D6434FF9417456C113B2B59750EE [I3EC5B1B4C96DB2313F610F9A4300E221 ]; else
if (I9ED39E2EA931586B6A985A6942EF573E == I5C62905D226C50178205CCCDB8C82788 ) begin if (I93707F725009F066ECF17DD8F6409A66 ) IE9E97C511899C07C74E75269A2ABA956
= 8'b101_11100; else IE9E97C511899C07C74E75269A2ABA956 = IC253D6434FF9417456C113B2B59750EE [I3EC5B1B4C96DB2313F610F9A4300E221 ]; end else
IE9E97C511899C07C74E75269A2ABA956 = 8'b001_11100; end always @(*) begin if ( I9ED39E2EA931586B6A985A6942EF573E ==
IE44F9E348E41CB272EFA87387728571B || (I9ED39E2EA931586B6A985A6942EF573E == I5C62905D226C50178205CCCDB8C82788 &&
!I93707F725009F066ECF17DD8F6409A66 ) ) begin I10315042C15E5BE9C16B02711AC72209 = 0; IB9C5339A9F988BDA02C82F2B8C804151
= IC253D6434FF9417456C113B2B59750EE [I3EC5B1B4C96DB2313F610F9A4300E221 ]; end else begin I10315042C15E5BE9C16B02711AC72209
= 1; IB9C5339A9F988BDA02C82F2B8C804151 = IA55086E1186D1C3CC0FFF510278DF91E ; end end logic [2:0] IB71403807C90F49A005DED2EC690370F ; always
@(posedge ID5972F1602659028768AC47B9316B673 ) if (I86266EE937D97F812A8E57D22B62EE29 ) IB71403807C90F49A005DED2EC690370F
<= {3{2'b00}}; else IB71403807C90F49A005DED2EC690370F <= {3{I363515199821A877761C5143490995BD }}; assign I021CFCAE834FA766B3091B6B708D8140
= ( ( IB71403807C90F49A005DED2EC690370F [0] & IB71403807C90F49A005DED2EC690370F [1] ) | ( IB71403807C90F49A005DED2EC690370F [1]
& IB71403807C90F49A005DED2EC690370F [2] ) | ( IB71403807C90F49A005DED2EC690370F [0] & IB71403807C90F49A005DED2EC690370F [2]
) ); logic [9:0] I3B1EDBF79F19D4A39E09A4A5BE990693 ; IABC6B35F4B0413305137538EE4407E67 I363BDF953355168947BD8B3FBF691BC0 (
.I02F62FEAFD6D93D552D5B8716C48A42B (IE9E97C511899C07C74E75269A2ABA956 ), .I8CE4B16B22B58894AA86C421E8759DF3 (I10315042C15E5BE9C16B02711AC72209 ),
.I1816A803A42A3A548A47FD7B90407CAC (I021CFCAE834FA766B3091B6B708D8140 ), .I8F9C634FB2FBC4B39107A845EF6445C6 (I3B1EDBF79F19D4A39E09A4A5BE990693 ),
.I8CD2DE889F491A5FFB5BB3AF153546D5 (I363515199821A877761C5143490995BD )); logic IEC4D1EB36B22D19728E9D1D23CA84D1C ; logic
[9:0] IA19F9F3EB524F6474AD00F1C2553C963 ; integer I865C0C0B4AB0E063E5CAA3387C1A8741 ; always @(*) begin case (IAD05C732EFA7E73CEB25AFAF7B6B2684 )
1'b0 : begin IA19F9F3EB524F6474AD00F1C2553C963 = {IB9C5339A9F988BDA02C82F2B8C804151 , 2'b0}; end 1'b1 : begin for
(I865C0C0B4AB0E063E5CAA3387C1A8741 =0; I865C0C0B4AB0E063E5CAA3387C1A8741 <10; I865C0C0B4AB0E063E5CAA3387C1A8741 =I865C0C0B4AB0E063E5CAA3387C1A8741 +1) IA19F9F3EB524F6474AD00F1C2553C963 [(10-1)-I865C0C0B4AB0E063E5CAA3387C1A8741 ]
= I3B1EDBF79F19D4A39E09A4A5BE990693 [I865C0C0B4AB0E063E5CAA3387C1A8741 ]; end endcase end logic I189154CAE37F6F62B37160F49AFB83C5 ,
I72B2B9DA666B665EA9F6986E481E852E ; assign I189154CAE37F6F62B37160F49AFB83C5 = I0A3BC2148686F2B562665C3891507E35 ;
assign ID5972F1602659028768AC47B9316B673 = I72B2B9DA666B665EA9F6986E481E852E ; logic [9:0] I780C2AA6563151EFA2CB302AA0DB9639 ; always @(posedge
ID5972F1602659028768AC47B9316B673 ) I780C2AA6563151EFA2CB302AA0DB9639 <= IA19F9F3EB524F6474AD00F1C2553C963 ; wire
I2C1D866ED67626BD73A37A83281336C8 ; I39607C0DCC66F95CC21E6ACF9889D96F I69897239BF3436DAD8887FDC9D29B69F (.I0A3BC2148686F2B562665C3891507E35 (I189154CAE37F6F62B37160F49AFB83C5 )
, .IF927D8348D0B86E1E1452C2EEF729055 (IAD05C732EFA7E73CEB25AFAF7B6B2684 ), .IC68271A63DDBC431C307BEB7D2918275 (I72B2B9DA666B665EA9F6986E481E852E ),
.IEC4D1EB36B22D19728E9D1D23CA84D1C (IEC4D1EB36B22D19728E9D1D23CA84D1C )); I84F6FB7CD5CD53B5679489A29396448F I4D5EF19F9F4836EB24F6EA49892B1084
(.I0A3BC2148686F2B562665C3891507E35 (I189154CAE37F6F62B37160F49AFB83C5 ), .IEC4D1EB36B22D19728E9D1D23CA84D1C (IEC4D1EB36B22D19728E9D1D23CA84D1C ),
.I13B5BFE96F3E2FE411C9F66F4A582ADF (I780C2AA6563151EFA2CB302AA0DB9639 ), .IC68271A63DDBC431C307BEB7D2918275 (I2C1D866ED67626BD73A37A83281336C8 )); always @(*)
begin case (IB4702C9059470087164094C2E5F94070 ) 1'b1: begin IC68271A63DDBC431C307BEB7D2918275 = I0A3BC2148686F2B562665C3891507E35 ;
end 1'b0: begin IC68271A63DDBC431C307BEB7D2918275 = I2C1D866ED67626BD73A37A83281336C8 ; end endcase end endmodule

